../../VGA/VGA_Vsync_gen.vhd