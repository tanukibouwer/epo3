configuration chip_toplevel_routed_cfg of chip_toplevel is
   for routed
      -- skipping del01bwp7t because it is not a local entity
      -- skipping ckbd0bwp7t because it is not a local entity
      -- skipping del1bwp7t because it is not a local entity
      -- skipping del0bwp7t because it is not a local entity
      -- skipping del02bwp7t because it is not a local entity
      -- skipping del2bwp7t because it is not a local entity
      -- skipping buffd1p5bwp7t because it is not a local entity
      -- skipping buffd2bwp7t because it is not a local entity
      -- skipping ckbd12bwp7t because it is not a local entity
      -- skipping ckbd8bwp7t because it is not a local entity
      -- skipping invd2bwp7t because it is not a local entity
      -- skipping invd1bwp7t because it is not a local entity
      -- skipping invd0bwp7t because it is not a local entity
      for all: orientation use configuration work.orientation_behavioural_cfg;
      end for;
      for all: input_period_counter use configuration work.input_period_counter_behavioural_cfg;
      end for;
      -- skipping iao21d0bwp7t because it is not a local entity
      -- skipping or4d1bwp7t because it is not a local entity
      -- skipping ind3d1bwp7t because it is not a local entity
      -- skipping ao22d0bwp7t because it is not a local entity
      -- skipping aoi22d0bwp7t because it is not a local entity
      -- skipping ao32d0bwp7t because it is not a local entity
      -- skipping nd2d1bwp7t because it is not a local entity
      -- skipping aoi31d0bwp7t because it is not a local entity
      -- skipping dfkcnqd1bwp7t because it is not a local entity
      -- skipping dfqd1bwp7t because it is not a local entity
      -- skipping edfkcnqd1bwp7t because it is not a local entity
      -- skipping ao221d0bwp7t because it is not a local entity
      -- skipping moai22d0bwp7t because it is not a local entity
      -- skipping ao211d0bwp7t because it is not a local entity
      -- skipping oai31d0bwp7t because it is not a local entity
      -- skipping oai21d0bwp7t because it is not a local entity
      -- skipping oa21d0bwp7t because it is not a local entity
      -- skipping nr3d0bwp7t because it is not a local entity
      -- skipping oai221d1bwp7t because it is not a local entity
      -- skipping oa211d0bwp7t because it is not a local entity
      -- skipping nd4d0bwp7t because it is not a local entity
      -- skipping oai211d1bwp7t because it is not a local entity
      -- skipping nr2xd0bwp7t because it is not a local entity
      -- skipping oai222d0bwp7t because it is not a local entity
      -- skipping aoi33d1bwp7t because it is not a local entity
      -- skipping aoi221d0bwp7t because it is not a local entity
      -- skipping aoi211xd0bwp7t because it is not a local entity
      -- skipping or3d1bwp7t because it is not a local entity
      -- skipping aoi21d0bwp7t because it is not a local entity
      -- skipping nr4d0bwp7t because it is not a local entity
      -- skipping nr2d1bwp7t because it is not a local entity
      -- skipping maoi22d0bwp7t because it is not a local entity
      -- skipping or2d1bwp7t because it is not a local entity
      -- skipping ao21d0bwp7t because it is not a local entity
      -- skipping maoi222d1bwp7t because it is not a local entity
      -- skipping nd3d0bwp7t because it is not a local entity
      -- skipping inr3d0bwp7t because it is not a local entity
      -- skipping ckxor2d1bwp7t because it is not a local entity
      -- skipping fa1d0bwp7t because it is not a local entity
      -- skipping ind2d1bwp7t because it is not a local entity
      -- skipping inr2d1bwp7t because it is not a local entity
      -- skipping oai22d0bwp7t because it is not a local entity
      -- skipping oai221d0bwp7t because it is not a local entity
      -- skipping oai31d1bwp7t because it is not a local entity
      -- skipping nr2d0bwp7t because it is not a local entity
      -- skipping an2d0bwp7t because it is not a local entity
      -- skipping ha1d0bwp7t because it is not a local entity
      -- skipping aoi211d0bwp7t because it is not a local entity
      -- skipping inr2xd0bwp7t because it is not a local entity
      -- skipping inr2d0bwp7t because it is not a local entity
      -- skipping cknd1bwp7t because it is not a local entity
      -- skipping aoi222d0bwp7t because it is not a local entity
      -- skipping an4d0bwp7t because it is not a local entity
      -- skipping ckmux2d1bwp7t because it is not a local entity
      -- skipping ioa21d0bwp7t because it is not a local entity
      -- skipping xnr2d1bwp7t because it is not a local entity
      -- skipping nr2d1p5bwp7t because it is not a local entity
      -- skipping nd4d1bwp7t because it is not a local entity
      -- skipping nd2d0bwp7t because it is not a local entity
      -- skipping an2d1bwp7t because it is not a local entity
      -- skipping iinr4d0bwp7t because it is not a local entity
      -- skipping oa22d0bwp7t because it is not a local entity
      -- skipping dfd1bwp7t because it is not a local entity
      -- skipping ao31d1bwp7t because it is not a local entity
      -- skipping cknd2d1bwp7t because it is not a local entity
      -- skipping xor3d1bwp7t because it is not a local entity
      -- skipping ind4d0bwp7t because it is not a local entity
      -- skipping oa32d1bwp7t because it is not a local entity
      -- skipping aoi221d1bwp7t because it is not a local entity
      -- skipping an3d1bwp7t because it is not a local entity
      -- skipping an3d0bwp7t because it is not a local entity
      -- skipping inr4d0bwp7t because it is not a local entity
      -- skipping oa221d0bwp7t because it is not a local entity
      -- skipping ioa21d1bwp7t because it is not a local entity
      -- skipping oa222d0bwp7t because it is not a local entity
      -- skipping oai32d1bwp7t because it is not a local entity
      -- skipping oai32d0bwp7t because it is not a local entity
      -- skipping oa33d0bwp7t because it is not a local entity
      -- skipping ind3d0bwp7t because it is not a local entity
      -- skipping ckan2d1bwp7t because it is not a local entity
      -- skipping xor4d1bwp7t because it is not a local entity
      -- skipping ao32d1bwp7t because it is not a local entity
      -- skipping ao222d0bwp7t because it is not a local entity
      -- skipping aoi32d1bwp7t because it is not a local entity
      -- skipping dfkcnd1bwp7t because it is not a local entity
      -- skipping invd5bwp7t because it is not a local entity
      -- skipping dfqd0bwp7t because it is not a local entity
      -- skipping ckan2d8bwp7t because it is not a local entity
      -- skipping oa31d1bwp7t because it is not a local entity
      -- skipping edfkcnd1bwp7t because it is not a local entity
      -- skipping dfksnd1bwp7t because it is not a local entity
      -- skipping an4d1bwp7t because it is not a local entity
      -- skipping dfd0bwp7t because it is not a local entity
      -- skipping cknd10bwp7t because it is not a local entity
      -- skipping aoi211d1bwp7t because it is not a local entity
      -- skipping oai33d1bwp7t because it is not a local entity
      -- skipping ind2d0bwp7t because it is not a local entity
      -- skipping nd3d1bwp7t because it is not a local entity
      -- skipping or4xd1bwp7t because it is not a local entity
      -- skipping aoi21d1bwp7t because it is not a local entity
      -- skipping iind4d0bwp7t because it is not a local entity
      -- skipping dfxd1bwp7t because it is not a local entity
      -- skipping ind4d1bwp7t because it is not a local entity
   end for;
end chip_toplevel_routed_cfg;
