../../attack/attackpressed-behavioural-cfg.vhd