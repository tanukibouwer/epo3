../../memory/m_ram4bit_cfg.vhd