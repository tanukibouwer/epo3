--module: char_sprite
--version: 1
--author: Parama Fawwaz 
--------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------
--MODULE DESCRIPTION
--! This module is the static ROM for the sprites regarding the character frames that can be shown on screen
--! 
--! This will be a modular component with an enable signal that will allow for the component to take over
--! coloring duties
--! 
--------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity char_sprites is
    port (
        reset  : in std_logic;
        sprite: in std_logic_vector(3 downto 0); -- 9 (max is 1001 in binary)
        


        R_data : out std_logic_vector(3 downto 0);
        G_data : out std_logic_vector(3 downto 0);
        B_data : out std_logic_vector(3 downto 0)

    );
end char_sprites;

--table:
-- sprite = 0: jump/crouch sprite
-- sprite = 1: running sprite 1
-- sprite = 2: running sprite 2
-- sprite = 3: running sprite 3


architecture behavioural of char_sprites is

    -- declare the array for the colours --> copy from number_sprite.vhd basically, but different sprites
    subtype color_val is std_logic_vector(11 downto 0); -- R(11,10,9,8) G(7,6,5,4) B(3,2,1,0)
    type char_sprite_x is array (0 to 7) of color_val;
    type char_sprite_y is array (0 to 11) of char_sprite_x;

    -- fill the arrays
    constant zero : char_sprite_y := ( 
        (("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011")), 
        (("001101100011"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
        (("001101100011"),("111111111111"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011")), 
        (("001101100011"),("111111111111"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011")), 
        (("001101100011"),("111111111111"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011")), 
        (("001101100011"),("111111111111"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011")), 
        (("001101100011"),("111111111111"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011")), 
        (("001101100011"),("111111111111"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011")), 
        (("001101100011"),("111111111111"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011")), 
        (("001101100011"),("111111111111"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011")),         
        (("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011"),("001101100011")) 
    ); 

    constant running_1 : char_sprite_y := (
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("110000100001"),("110000100001"),("110000100001"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("110000100001"),("110000100001"),("110000100001"),("110000100001")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("111111111111"),("111111111111"),("000000000000"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("111111111111"),("111111111111"),("000000000000"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("111111111111"),("111111111111"),("111111111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("110000100001"),("110000100001"),("110000100001"),("000010111111"),("000010111111"),("111111111111")),
        (
        ("000010111111"),("110000100001"),("000010111111"),("110000100001"),("110000100001"),("110000100001"),("110000100001"),("000010111111")),
        (
        ("111111111111"),("000010111111"),("000010111111"),("110000100001"),("110000100001"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("110000100001"),("110000100001"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("110000100001"),("000010111111"),("110000100001"),("110000100001"),("000010111111"),("000010111111")),
        (
        ("111111111111"),("110000100001"),("000010111111"),("000010111111"),("000010111111"),("000010111111"),("110000100001"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111"),("111111111111"),("000010111111"))
        )
    begin 
    case sprite is
        when "0001"

end behavioural;