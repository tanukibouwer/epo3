configuration attackpressed_behavioural_cfg of attackp is
	for behavioural
		end for;
end configuration attackpressed_behavioural_cfg;
