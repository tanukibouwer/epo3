configuration coloring_cfg of coloring is
    for structural
    end for;
end configuration coloring_cfg;