../../physics/collision_resolver.vhd