../../physics/h_player_movement_behaviour_cfg.vhd