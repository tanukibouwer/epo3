configuration char_animation_fsm_cfg of char_animation_fsm is
    for behavioural
        for all : frame_cnt use work.frame_cnt_cfg; 
    end for;
end configuration char_animation_fsm_cfg;