configuration V_line_cnt_cfg of v_line_cnt is
    for behavioural
    end for;
end configuration V_line_cnt_cfg;