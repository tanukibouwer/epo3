../../physics/position_adder_behaviour_cfg.vhd