configuration physics_system_tb_behaviour_cfg of physics_system_tb is
   for behaviour
      for all: physics_system use configuration work.physics_system_behaviour_cfg;
      end for;
   end for;
end physics_system_tb_behaviour_cfg;
