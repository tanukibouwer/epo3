configuration collision_resolver_behaviour_cfg of collision_resolver is
   for behaviour
   end for;
end collision_resolver_behaviour_cfg;
