../../attack/damagecalculator-behavioural-cfg.vhd