../../attack/orientation-behavioural-cfg.vhd