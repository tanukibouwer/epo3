--module: char_sprite
--version: 1
--author: Parama Fawwaz & Kevin Vermaat
--------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------
--MODULE DESCRIPTION
--! This module is the static ROM for the sprites regarding the character frames that can be shown on screen
--! 
--! This will be a modular component with an enable signal that will allow for the component to take over
--! coloring duties
--! 
-- 
-- Notes:
-- for the controller inputs, take note of the following
-- bit 3 is down, bit 2 is jump, bit 1 is right, bit 0 is left
-- others are as of now not required
--------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity char_sprites is
    port (
        -- global or constant control signals
        clk   : in std_logic;
        reset : in std_logic;
        player : in std_logic; 
        -- controller input information
        orientation : in std_logic;
        controller  : in std_logic_vector(7 downto 0);
        -- going through the array
        -- count for where one is
        hcount : in std_logic_vector(9 downto 0);
        vcount : in std_logic_vector(9 downto 0);
        -- top and left bounds for normalisation
        boundx : in std_logic_vector(9 downto 0);
        boundy : in std_logic_vector(9 downto 0);

        -- RGB outputs
        R_data : out std_logic_vector(3 downto 0);
        G_data : out std_logic_vector(3 downto 0);
        B_data : out std_logic_vector(3 downto 0)

    );
end char_sprites;
architecture behavioural of char_sprites is

    component char_animation_fsm is
        port (
            clk   : in std_logic;
            reset : in std_logic;

            -- global frame counters
            vcount : in std_logic_vector(9 downto 0); -- vertical frame counter
            hcount : in std_logic_vector(9 downto 0); -- horizontal line counter

            -- controller input signal
            controller_in : in std_logic_vector(7 downto 0); -- bit 0 = left, bit 1 = right, bit 2 = up, bit 3 = down

            -- sprite output value
            sprite : out std_logic_vector(1 downto 0)
        );
    end component;

    -- control signals for the animation fsm
    -- signal an_on  : std_logic;
    -- signal frame  : std_logic;
    signal sprite : std_logic_vector(1 downto 0);

    -- integer values for the counts
    -- signal int_hcount, int_vcount : integer;
    -- signal int_boundx, int_boundy : integer;

    -- declare the array for the colours --> copy from number_sprite.vhd basically, but different sprites --> for now sprite left and right is the same for now
    constant sprite_x_length : integer := 31;
    constant sprite_y_length : integer := 47;
    subtype color_val is std_logic_vector(11 downto 0); -- R(11,10,9,8) G(7,6,5,4) B(3,2,1,0)
    type char_sprite_x is array (0 to sprite_x_length) of color_val;
    type char_sprite_y is array (0 to sprite_y_length) of char_sprite_x;

    -- fill the arrays
    constant running_1 : char_sprite_y :=
        ( 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("000000000000"),("000000000000"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("000000000000"),("000000000000"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("101110111011"),("101110111011"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("111111101100"),("111111101100"),("111111101100")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("111111101100"),("111111101100"),("111111101100")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("111111101100"),("111111101100"),("111111101100")), 
        (("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("111111101100"),("111111101100"),("111111101100")), 
        (("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111")), 
        (("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111")), 
        (("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111")), 
        (("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111")), 
        (("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111")), 
        (("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111")), 
        (("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111")), 
        (("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001")) 
    ); 
    constant idle_1 : char_sprite_y := 
        ( 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("000000000000"),("000000000000"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("000000000000"),("000000000000"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("101110111011"),("101110111011"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("111011011011"),("111011011011"),("111011011011"),("111011011011"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("111011011011"),("111011011011"),("111011011011"),("111011011011"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("111011011011"),("111011011011"),("111011011011"),("111011011011"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("111011011011"),("111011011011"),("111011011011"),("111011011011"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")) 
    ); 
    constant jump_crouch_1 : char_sprite_y := 
        ( 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("000000000000"),("000000000000"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("000000000000"),("000000000000"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("101110111011"),("101110111011"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("111011011011"),("111011011011"),("111011011011"),("111011011011"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("111011011011"),("111011011011"),("111011011011"),("111011011011"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("111011011011"),("111011011011"),("111011011011"),("111011011011"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("111011011011"),("111011011011"),("111011011011"),("111011011011"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("111011011011"),("111011011011"),("111011011011"),("111011011011"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("111011011011"),("111011011011"),("111011011011"),("111011011011"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("111011011011"),("111011011011"),("111011011011"),("111011011011"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("111011011011"),("111011011011"),("111011011011"),("111011011011"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")) 
    ); 
    constant running_2 : char_sprite_y := 
        ( 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("111011010110"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000000000000"),("000000000000"),("111111111111"),("111111111111"),("111111101100"),("111011010110"),("111011010110"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000000000000"),("000000000000"),("111111111111"),("111111111111"),("111111101100"),("111011010110"),("111011010110"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000000000000"),("000000000000"),("111111111111"),("111111111111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000000000000"),("000000000000"),("111111111111"),("111111111111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100")), 
        (("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100")), 
        (("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100")), 
        (("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100")), 
        (("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100")), 
        (("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100")), 
        (("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100")) 
    ); 
    constant idle_2 : char_sprite_y := 
        ( 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("111011010110"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000000000000"),("000000000000"),("111111111111"),("111111111111"),("111111101100"),("111011010110"),("111011010110"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000000000000"),("000000000000"),("111111111111"),("111111111111"),("111111101100"),("111011010110"),("111011010110"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000000000000"),("000000000000"),("111111111111"),("111111111111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000000000000"),("000000000000"),("111111111111"),("111111111111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")) 
    ); 
    constant jump_crouch_2 : char_sprite_y := 
        ( 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("111011010110"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000000000000"),("000000000000"),("111111111111"),("111111111111"),("111111101100"),("111011010110"),("111011010110"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000000000000"),("000000000000"),("111111111111"),("111111111111"),("111111101100"),("111011010110"),("111011010110"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000000000000"),("000000000000"),("111111111111"),("111111111111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000000000000"),("000000000000"),("111111111111"),("111111111111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")) 
    ); 
    constant attack_1 : char_sprite_y := ( 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("101010101010"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("000000000000"),("000000000000"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("101010101010"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("000000000000"),("000000000000"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("101110111011"),("101110111011"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("111111101100"),("111111101100"),("111111101100"),("111111101100")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("111111101100"),("111111101100"),("111111101100"),("111111101100")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("111111101100"),("111111101100"),("111111101100"),("111111101100")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("111111101100"),("111111101100"),("111111101100"),("111111101100")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("011001010101"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("011110011001"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")) 
    ); 
    constant attack_2 : char_sprite_y :=( 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("111011010110"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000000000000"),("000000000000"),("111111111111"),("111111111111"),("111111101100"),("111011010110"),("111011010110"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000000000000"),("000000000000"),("111111111111"),("111111111111"),("111111101100"),("111011010110"),("111011010110"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000000000000"),("000000000000"),("111111111111"),("111111111111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000000000000"),("000000000000"),("111111111111"),("111111111111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111011010110"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("111111101100"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("111111101100"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("111111101100"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("111111101100"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("111111101100"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("111111101100"),("111111101100"),("111111101100"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("011110010111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")), 
        (("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("011101010100"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111"),("000011001111")) 
    ); 
begin
    -- int_hcount <= to_integer(unsigned(hcount));
    -- int_vcount <= to_integer(unsigned(vcount));
    -- int_boundx <= to_integer(unsigned(boundx));
    -- int_boundy <= to_integer(unsigned(boundy));

    frame_control : char_animation_fsm port map(
        clk           => clk,
        reset         => reset,
        vcount        => vcount,
        hcount        => hcount,
        controller_in => controller,
        sprite        => sprite
    );

    process (sprite, orientation, player, hcount, vcount, boundx, boundy)
        variable int_boundx : integer;
        variable int_boundy : integer;
        variable int_hcount : integer;
        variable int_vcount : integer;
    begin
        int_hcount := to_integer(unsigned(hcount));
        int_vcount := to_integer(unsigned(vcount));
        int_boundx := to_integer(unsigned(boundx));
        int_boundy := to_integer(unsigned(boundy));

        -- choose which "animation" to play dependent on the input
        -- R_data <= jump_crouch_R(int_vcount - (int_boundy))(int_hcount - (int_boundx))(11 downto 8);
        -- G_data <= jump_crouch_R(int_vcount - (int_boundy))(int_hcount - (int_boundx))(7 downto 4);
        -- B_data <= jump_crouch_R(int_vcount - (int_boundy))(int_hcount - (int_boundx))(3 downto 0);
        case sprite is
            when "00" => -- show idle sprite
                if orientation = '1' then -- show the sprite how it is drawn
                    if player = '0' then -- if it is player 1 then show the sprite for player 2
                        R_data <= idle_1(int_vcount - (int_boundy))(int_hcount - (int_boundx))(11 downto 8);
                        G_data <= idle_1(int_vcount - (int_boundy))(int_hcount - (int_boundx))(7 downto 4);
                        B_data <= idle_1(int_vcount - (int_boundy))(int_hcount - (int_boundx))(3 downto 0);
                    else --  if it is player 2 then show the sprite for player 2
                        R_data <= idle_2(int_vcount - (int_boundy))(sprite_x_length - (int_hcount - (int_boundx)))(11 downto 8);
                        G_data <= idle_2(int_vcount - (int_boundy))(sprite_x_length - (int_hcount - (int_boundx)))(7 downto 4);
                        B_data <= idle_2(int_vcount - (int_boundy))(sprite_x_length - (int_hcount - (int_boundx)))(3 downto 0);
                    end if;
                elsif orientation = '0' then -- show the sprite in verted to how it is drawn
                    if player = '0' then -- if it is player 1 then show the sprite for player 2
                        R_data <= idle_1((int_vcount - (int_boundy)))(sprite_x_length - (int_hcount - (int_boundx)))(11 downto 8);
                        G_data <= idle_1((int_vcount - (int_boundy)))(sprite_x_length - (int_hcount - (int_boundx)))(7 downto 4);
                        B_data <= idle_1((int_vcount - (int_boundy)))(sprite_x_length - (int_hcount - (int_boundx)))(3 downto 0);
                    else --  if it is player 2 then show the sprite for player 2
                        R_data <= idle_2((int_vcount - (int_boundy)))(int_hcount - (int_boundx))(11 downto 8);
                        G_data <= idle_2((int_vcount - (int_boundy)))(int_hcount - (int_boundx))(7 downto 4);
                        B_data <= idle_2((int_vcount - (int_boundy)))(int_hcount - (int_boundx))(3 downto 0);
                    end if;
                else 
                    R_data <= "0000";
                    G_data <= "0000";
                    B_data <= "0000";    
                end if;
            when "01" => -- show ducking sprite
                if orientation = '1' then -- show the sprite how it is drawn
                    if player = '0' then -- if it is player 1 then show the sprite for player 2
                        R_data <= jump_crouch_1(int_vcount - (int_boundy))(int_hcount - (int_boundx))(11 downto 8);
                        G_data <= jump_crouch_1(int_vcount - (int_boundy))(int_hcount - (int_boundx))(7 downto 4);
                        B_data <= jump_crouch_1(int_vcount - (int_boundy))(int_hcount - (int_boundx))(3 downto 0);
                    else --  if it is player 2 then show the sprite for player 2
                        R_data <= jump_crouch_2(int_vcount - (int_boundy))(sprite_x_length - (int_hcount - (int_boundx)))(11 downto 8);
                        G_data <= jump_crouch_2(int_vcount - (int_boundy))(sprite_x_length - (int_hcount - (int_boundx)))(7 downto 4);
                        B_data <= jump_crouch_2(int_vcount - (int_boundy))(sprite_x_length - (int_hcount - (int_boundx)))(3 downto 0);
                    end if;
                elsif orientation = '0' then -- show the sprite in verted to how it is drawn
                    if player = '0' then -- if it is player 1 then show the sprite for player 2
                        R_data <= jump_crouch_1((int_vcount - (int_boundy)))(sprite_x_length - (int_hcount - (int_boundx)))(11 downto 8);
                        G_data <= jump_crouch_1((int_vcount - (int_boundy)))(sprite_x_length - (int_hcount - (int_boundx)))(7 downto 4);
                        B_data <= jump_crouch_1((int_vcount - (int_boundy)))(sprite_x_length - (int_hcount - (int_boundx)))(3 downto 0);
                    else --  if it is player 2 then show the sprite for player 2
                        R_data <= jump_crouch_2((int_vcount - (int_boundy)))(int_hcount - (int_boundx))(11 downto 8);
                        G_data <= jump_crouch_2((int_vcount - (int_boundy)))(int_hcount - (int_boundx))(7 downto 4);
                        B_data <= jump_crouch_2((int_vcount - (int_boundy)))(int_hcount - (int_boundx))(3 downto 0);
                    end if;
                else 
                    R_data <= "0000";
                    G_data <= "0000";
                    B_data <= "0000";    
                end if;
            when "10" => -- show running sprite
                if orientation = '1' then -- show the sprite how it is drawn
                    if player = '0' then -- if it is player 1 then show the sprite for player 2
                        R_data <= running_1(int_vcount - (int_boundy))(int_hcount - (int_boundx))(11 downto 8);
                        G_data <= running_1(int_vcount - (int_boundy))(int_hcount - (int_boundx))(7 downto 4);
                        B_data <= running_1(int_vcount - (int_boundy))(int_hcount - (int_boundx))(3 downto 0);
                    else --  if it is player 2 then show the sprite for player 2
                        R_data <= running_2(int_vcount - (int_boundy))(sprite_x_length - (int_hcount - (int_boundx)))(11 downto 8);
                        G_data <= running_2(int_vcount - (int_boundy))(sprite_x_length - (int_hcount - (int_boundx)))(7 downto 4);
                        B_data <= running_2(int_vcount - (int_boundy))(sprite_x_length - (int_hcount - (int_boundx)))(3 downto 0);
                    end if;
                elsif orientation = '0' then -- show the sprite in verted to how it is drawn
                    if player = '0' then -- if it is player 1 then show the sprite for player 2
                        R_data <= running_1((int_vcount - (int_boundy)))(sprite_x_length - (int_hcount - (int_boundx)))(11 downto 8);
                        G_data <= running_1((int_vcount - (int_boundy)))(sprite_x_length - (int_hcount - (int_boundx)))(7 downto 4);
                        B_data <= running_1((int_vcount - (int_boundy)))(sprite_x_length - (int_hcount - (int_boundx)))(3 downto 0);
                    else --  if it is player 2 then show the sprite for player 2
                        R_data <= running_2((int_vcount - (int_boundy)))(int_hcount - (int_boundx))(11 downto 8);
                        G_data <= running_2((int_vcount - (int_boundy)))(int_hcount - (int_boundx))(7 downto 4);
                        B_data <= running_2((int_vcount - (int_boundy)))(int_hcount - (int_boundx))(3 downto 0);
                    end if;
                else 
                    R_data <= "0000";
                    G_data <= "0000";
                    B_data <= "0000";    
                end if;
            when "11" => 
            if orientation = '1' then -- show the sprite how it is drawn
                if player = '0' then -- if it is player 1 then show the sprite for player 2
                    R_data <= attack_1(int_vcount - (int_boundy))(int_hcount - (int_boundx))(11 downto 8);
                    G_data <= attack_1(int_vcount - (int_boundy))(int_hcount - (int_boundx))(7 downto 4);
                    B_data <= attack_1(int_vcount - (int_boundy))(int_hcount - (int_boundx))(3 downto 0);
                else --  if it is player 2 then show the sprite for player 2
                    R_data <= attack_2(int_vcount - (int_boundy))(sprite_x_length - (int_hcount - (int_boundx)))(11 downto 8);
                    G_data <= attack_2(int_vcount - (int_boundy))(sprite_x_length - (int_hcount - (int_boundx)))(7 downto 4);
                    B_data <= attack_2(int_vcount - (int_boundy))(sprite_x_length - (int_hcount - (int_boundx)))(3 downto 0);
                end if;
            elsif orientation = '0' then -- show the sprite in verted to how it is drawn
                if player = '0' then -- if it is player 1 then show the sprite for player 2
                    R_data <= attack_1((int_vcount - (int_boundy)))(sprite_x_length - (int_hcount - (int_boundx)))(11 downto 8);
                    G_data <= attack_1((int_vcount - (int_boundy)))(sprite_x_length - (int_hcount - (int_boundx)))(7 downto 4);
                    B_data <= attack_1((int_vcount - (int_boundy)))(sprite_x_length - (int_hcount - (int_boundx)))(3 downto 0);
                else --  if it is player 2 then show the sprite for player 2
                    R_data <= attack_2((int_vcount - (int_boundy)))(int_hcount - (int_boundx))(11 downto 8);
                    G_data <= attack_2((int_vcount - (int_boundy)))(int_hcount - (int_boundx))(7 downto 4);
                    B_data <= attack_2((int_vcount - (int_boundy)))(int_hcount - (int_boundx))(3 downto 0);
                end if;
            else 
                R_data <= "0000";
                G_data <= "0000";
                B_data <= "0000";    
            end if;

            when others =>
                R_data <= "0000";
                G_data <= "0000";
                B_data <= "0000";

        end case;
    end process;

end behavioural;