configuration gravity_tb_structural_cfg of gravity_tb is
   for structural
      for all: gravity use configuration work.gravity_behaviour_cfg;
      end for;
   end for;
end gravity_tb_structural_cfg;
