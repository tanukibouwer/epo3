../../VGA/VGA_number_sprite.vhd