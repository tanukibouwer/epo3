configuration input_deserializer_behavioural_cfg of input_deserializer is
	for behavioural
		end for;
end configuration input_deserializer_behavioural_cfg;
