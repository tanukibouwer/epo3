../../memory/m_ram10bit.vhd