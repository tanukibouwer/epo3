../../input/input_register_behavioural_cfg.vhd