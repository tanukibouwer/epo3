--module: char_sprite
--version: 1
--author: Parama Fawwaz 
--------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------
--MODULE DESCRIPTION
--! This module is the static ROM for the sprites regarding the character frames that can be shown on screen
--! 
--! This will be a modular component with an enable signal that will allow for the component to take over
--! coloring duties
--! 
--------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity char_sprites is
    port (
        reset  : in std_logic;
        sprite: in std_logic_vector(2 downto 0); -- 9 (max is 1001 in binary)

        hcount : in std_logic_vector(9 downto 0);
        vcount : in std_logic_vector(9 downto 0);
        boundx : in std_logic_vector(9 downto 0);
        boundy : in std_logic_vector(9 downto 0);
        


        R_data : out std_logic_vector(3 downto 0);
        G_data : out std_logic_vector(3 downto 0);
        B_data : out std_logic_vector(3 downto 0)

    );
end char_sprites;


architecture behavioural of char_sprites is

    -- integer values for the counts
    signal int_hcount, int_vcount : integer;
    signal int_boundx, int_boundy : integer;

    -- declare the array for the colours --> copy from number_sprite.vhd basically, but different sprites
    subtype color_val is std_logic_vector(11 downto 0); -- R(11,10,9,8) G(7,6,5,4) B(3,2,1,0)
    type char_sprite_x is array (0 to 7) of color_val;
    type char_sprite_y is array (0 to 11) of char_sprite_x;

    -- fill the arrays
    constant running_1_R : char_sprite_y := (
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("110000010001"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("110000010001"),("110000010001")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("111111111111"),("111111111111"),("000000000000"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("111111111111"),("111111111111"),("000000000000"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("111111111111"),("111111111111"),("111111111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("110000010001"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("111111111111")),
        (
        ("000010111111"),("110000010001"),("000010111111"),("110000010001"),("110000010001"),("110000010001"),("110000010001"),("000010111111")),
        (
        ("111111111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("110000010001"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("000010111111")),
        (
        ("111111111111"),("110000010001"),("000010111111"),("000010111111"),("000010111111"),("000010111111"),("110000010001"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111"),("111111111111"),("000010111111"))
        );
    
    constant running_1_L : char_sprite_y := (
        (
        ("000010111111"),("110000010001"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("110000010001"),("110000010001"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000000000000"),("111111111111"),("111111111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000000000000"),("111111111111"),("111111111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("111111111111"),("111111111111"),("111111111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("111111111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("110000010001"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("110000010001"),("110000010001"),("110000010001"),("110000010001"),("000010111111"),("110000010001"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("111111111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("110000010001"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("110000010001"),("000010111111"),("000010111111"),("000010111111"),("000010111111"),("110000010001"),("111111111111")),
        (
        ("000010111111"),("111111111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111"))
        );

    constant idle_1_R : char_sprite_y := (
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("110000010001"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("110000010001"),("110000010001")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("111111111111"),("111111111111"),("000000000000"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("111111111111"),("111111111111"),("000000000000"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("111111111111"),("111111111111"),("111111111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("111111111111"),("110000010001"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("111111111111"),("111111111111"),("000010111111"),("000010111111"),("000010111111"))
        );

    constant idle_1_L : char_sprite_y := (
        (
        ("000010111111"),("110000010001"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("110000010001"),("110000010001"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000000000000"),("111111111111"),("111111111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000000000000"),("111111111111"),("111111111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("111111111111"),("111111111111"),("111111111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("110000010001"),("111111111111"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("111111111111"),("111111111111"),("000010111111"),("000010111111"),("000010111111"))
        );

    constant jump_crouch_R : char_sprite_y := (
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("110000010001"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("110000010001"),("110000010001")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("111111111111"),("111111111111"),("111111111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("111111111111"),("111111111111"),("000000000000"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("111111111111"),("111111111111"),("000000000000"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("110000010001"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("110000010001"),("111111111111"),("110000010001"),("111111111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("110000010001"),("110000010001"),("110000010001"),("110000010001"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("110000010001"),("000010111111"),("000010111111"),("111111111111"),("000010111111"),("000010111111")),
        (
        ("000010111111"),("000010111111"),("111111111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111"))
        );

        constant jump_crouch_L : char_sprite_y := (
            (
            ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
            (
            ("000010111111"),("110000010001"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
            (
            ("110000010001"),("110000010001"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
            (
            ("000010111111"),("000000000000"),("111111111111"),("111111111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
            (
            ("000010111111"),("000000000000"),("111111111111"),("111111111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
            (
            ("000010111111"),("111111111111"),("111111111111"),("111111111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111")),
            (
            ("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("110000010001"),("000010111111"),("000010111111")),
            (
            ("000010111111"),("000010111111"),("111111111111"),("110000010001"),("111111111111"),("110000010001"),("000010111111"),("000010111111")),
            (
            ("000010111111"),("000010111111"),("000010111111"),("110000010001"),("110000010001"),("000010111111"),("000010111111"),("000010111111")),
            (
            ("000010111111"),("000010111111"),("110000010001"),("110000010001"),("110000010001"),("110000010001"),("000010111111"),("000010111111")),
            (
            ("000010111111"),("000010111111"),("111111111111"),("000010111111"),("000010111111"),("110000010001"),("000010111111"),("000010111111")),
            (
            ("000010111111"),("000010111111"),("000010111111"),("000010111111"),("000010111111"),("111111111111"),("000010111111"),("000010111111"))
            );
    
--table:
-- sprite = 0: jump/crouch sprite right
-- sprite = 1: idle sprite 1 right
-- sprite = 2: running sprite 1 right
-- sprite = 3: jump/crouch sprite left
-- sprite = 4: idle sprite 1 left
-- sprite = 5: running sprite 1 left


begin 
    int_hcount <= to_integer(unsigned(hcount));
    int_vcount <= to_integer(unsigned(vcount));
    int_boundx <= to_integer(unsigned(boundx)) + 1;
    int_boundy <= to_integer(unsigned(boundy)) + 1;

    process (sprite, int_hcount, int_vcount, int_boundx, int_boundy)
    begin
        case sprite is
            when "000" => -- jump/crouch R
                R_data <= jump_crouch_R(int_vcount - int_boundy)(int_hcount - int_boundx)(11 downto 8);
                G_data <= jump_crouch_R(int_vcount - int_boundy)(int_hcount - int_boundx)(7 downto 4);
                B_data <= jump_crouch_R(int_vcount - int_boundy)(int_hcount - int_boundx)(3 downto 0);
            when "001" => -- idle1 R
                R_data <= idle_1_R(int_vcount - int_boundy)(int_hcount - int_boundx)(11 downto 8);
                G_data <= idle_1_R(int_vcount - int_boundy)(int_hcount - int_boundx)(7 downto 4);
                B_data <= idle_1_R(int_vcount - int_boundy)(int_hcount - int_boundx)(3 downto 0);
            when "010" => -- running1 R
                R_data <= running_1_R(int_vcount - int_boundy)(int_hcount - int_boundx)(11 downto 8);
                G_data <= running_1_R(int_vcount - int_boundy)(int_hcount - int_boundx)(7 downto 4);
                B_data <= running_1_R(int_vcount - int_boundy)(int_hcount - int_boundx)(3 downto 0);
            when "011" => -- jump/crouch L
                R_data <= jump_crouch_L(int_vcount - int_boundy)(int_hcount - int_boundx)(11 downto 8);
                G_data <= jump_crouch_L(int_vcount - int_boundy)(int_hcount - int_boundx)(7 downto 4);
                B_data <= jump_crouch_L(int_vcount - int_boundy)(int_hcount - int_boundx)(3 downto 0);
            when "100" => -- idle1 L
                R_data <= idle_1_L(int_vcount - int_boundy)(int_hcount - int_boundx)(11 downto 8);
                G_data <= idle_1_L(int_vcount - int_boundy)(int_hcount - int_boundx)(7 downto 4);
                B_data <= idle_1_L(int_vcount - int_boundy)(int_hcount - int_boundx)(3 downto 0);
            when "101" => -- running1 L
                R_data <= running_1_L(int_vcount - int_boundy)(int_hcount - int_boundx)(11 downto 8);
                G_data <= running_1_L(int_vcount - int_boundy)(int_hcount - int_boundx)(7 downto 4);
                B_data <= running_1_L(int_vcount - int_boundy)(int_hcount - int_boundx)(3 downto 0);

           
            when others => -- fallback for error handling and checking
                R_data <= "0000";
                G_data <= "0000";
                B_data <= "0000";
        end case;
    end process;

end behavioural;