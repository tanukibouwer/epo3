../../physics/gravity_behaviour_cfg.vhd