configuration hsync_gen_cfg of hsync_gen is
    for rtl
    end for;
end configuration hsync_gen_cfg;