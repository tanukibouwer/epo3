configuration number_sprite_cfg of number_sprite is
    for behavioural
    end for;
end configuration number_sprite_cfg;