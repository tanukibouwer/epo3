../../VGA/VGA_coloring_cfg.vhd