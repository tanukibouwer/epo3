configuration coldet_behaviour_cfg of coldet is
	for behaviour
	end for;
end configuraton coldet_behaviour_cfg;
