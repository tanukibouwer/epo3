configuration position_adder_behaviour_cfg of position_adder is
   for behaviour
   end for;
end position_adder_behaviour_cfg;
