../../VGA/VGA_dig3_num_splitter.vhd