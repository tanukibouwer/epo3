../../attack/coldet-behaviour.vhd