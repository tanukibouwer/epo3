../../VGA/VGA_Hsync_gen.vhd