../../main/t_8bregs.vhd