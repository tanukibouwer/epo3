--module: char_sprite
--version: 1
--author: Parama Fawwaz & Kevin Vermaat
--------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------
--MODULE DESCRIPTION
--! This module is the static ROM for the sprites regarding the character frames that can be shown on screen
--! 
--! This will be a modular component with an enable signal that will allow for the component to take over
--! coloring duties
--! 
-- 
-- Notes:
-- for the controller inputs, take note of the following
-- bit 3 is down, bit 2 is jump, bit 1 is right, bit 0 is left
-- others are as of now not required
--------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity char_sprites is
    port (
        clk   : in std_logic;
        reset : in std_logic;
        -- sprite control signals
        vsync_cnt   : in std_logic_vector(3 downto 0);
        orientation : in std_logic;
        controller  : in std_logic_vector(7 downto 0);
        -- going through the array
        hcount : in std_logic_vector(9 downto 0);
        vcount : in std_logic_vector(9 downto 0);
        boundx : in std_logic_vector(9 downto 0);
        boundy : in std_logic_vector(9 downto 0);

        R_data : out std_logic_vector(3 downto 0);
        G_data : out std_logic_vector(3 downto 0);
        B_data : out std_logic_vector(3 downto 0)

    );
end char_sprites;
architecture behavioural of char_sprites is

    component char_animation_fsm is
        port (
            clk   : in std_logic;
            reset : in std_logic;
            animation_clk : in std_logic_vector(3 downto 0);

            controller_in : in std_logic_vector(7 downto 0); -- bit 0 = left, bit 1 = right, bit 2 = up, bit 3 = down
            -- orientation   : in std_logic;                    --1 is right, 0 is left
            sprite : out std_logic_vector(1 downto 0)
            -- frame  : out std_logic
        );
    end component;

    -- control signals for the animation fsm
    signal an_on  : std_logic;
    -- signal frame  : std_logic;
    signal sprite : std_logic_vector(1 downto 0);

    -- integer values for the counts
    signal int_hcount, int_vcount : integer;
    signal int_boundx, int_boundy : integer;

    -- declare the array for the colours --> copy from number_sprite.vhd basically, but different sprites --> for now sprite left and right is the same for now
    subtype color_val is std_logic_vector(11 downto 0); -- R(11,10,9,8) G(7,6,5,4) B(3,2,1,0)
    type char_sprite_x is array (0 to 31) of color_val;
    type char_sprite_y is array (0 to 47) of char_sprite_x;

    -- fill the arrays
    constant running_1_R : char_sprite_y := (
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"))
    );
    constant running_1_L : char_sprite_y := (
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"))
    );
    constant idle_1_R : char_sprite_y := (
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"))
        );
        constant idle_1_L : char_sprite_y := (
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"))
    );
    constant jump_crouch_R : char_sprite_y := (
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"))
    );
    constant jump_crouch_L : char_sprite_y := (
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000000000000"), ("000000000000"), ("000000000000"), ("000000000000"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("110000010001"), ("110000010001"), ("110000010001"), ("110000010001"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111")),
        (
        ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("111111111111"), ("111111111111"), ("111111111111"), ("111111111111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"), ("000011001111"))
    );
    --table:
    -- sprite = 0: jump/crouch sprite right
    -- sprite = 1: idle sprite 1 right
    -- sprite = 2: running sprite 1 right
    -- sprite = 3: jump/crouch sprite left
    -- sprite = 4: idle sprite 1 left
    -- sprite = 5: running sprite 1 left
begin
    int_hcount <= to_integer(unsigned(hcount));
    int_vcount <= to_integer(unsigned(vcount));
    int_boundx <= to_integer(unsigned(boundx));
    int_boundy <= to_integer(unsigned(boundy));

    frame_control : char_animation_fsm port map(
        clk           => clk,
        reset         => reset,
        animation_clk => vsync_cnt,
        controller_in => controller,
        sprite        => sprite
    );

    process (sprite, orientation, int_hcount, int_vcount, int_boundx, int_boundy)
    begin
        -- choose which "animation" to play dependent on the input
        -- R_data <= jump_crouch_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(11 downto 8);
        -- G_data <= jump_crouch_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(7 downto 4);
        -- B_data <= jump_crouch_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(3 downto 0);
        case sprite is
            when "00" => -- show idle sprite
                if orientation = '0' then
                    R_data <= idle_1_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(11 downto 8);
                    G_data <= idle_1_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(7 downto 4);
                    B_data <= idle_1_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(3 downto 0);
                elsif orientation = '1' then
                    R_data <= idle_1_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(11 downto 8);
                    G_data <= idle_1_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(7 downto 4);
                    B_data <= idle_1_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(3 downto 0);
                end if;
            when "01" => -- show ducking sprite
                if orientation = '0' then
                    R_data <= jump_crouch_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(11 downto 8);
                    G_data <= jump_crouch_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(7 downto 4);
                    B_data <= jump_crouch_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(3 downto 0);
                elsif orientation = '1' then
                    R_data <= jump_crouch_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(11 downto 8);
                    G_data <= jump_crouch_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(7 downto 4);
                    B_data <= jump_crouch_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(3 downto 0);
                end if;
            when "10" => -- show running sprite
                if orientation = '0' then
                    R_data <= running_1_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(11 downto 8);
                    G_data <= running_1_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(7 downto 4);
                    B_data <= running_1_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(3 downto 0);
                elsif orientation = '1' then
                    R_data <= running_1_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(11 downto 8);
                    G_data <= running_1_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(7 downto 4);
                    B_data <= running_1_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(3 downto 0);
                end if;

            when others =>
                R_data <= "0000";
                G_data <= "0000";
                B_data <= "0000";

        end case;

        -- case vsync_cnt is
        --     when "000" => -- jump/crouch R
        --         R_data <= jump_crouch_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(11 downto 8);
        --         G_data <= jump_crouch_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(7 downto 4);
        --         B_data <= jump_crouch_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(3 downto 0);
        --     when "001" => -- idle1 R
        --         R_data <= idle_1_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(11 downto 8);
        --         G_data <= idle_1_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(7 downto 4);
        --         B_data <= idle_1_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(3 downto 0);
        --     when "010" => -- running1 R
        --         R_data <= running_1_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(11 downto 8);
        --         G_data <= running_1_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(7 downto 4);
        --         B_data <= running_1_R(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(3 downto 0);
        --     when "011" => -- jump/crouch L
        --         R_data <= jump_crouch_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(11 downto 8);
        --         G_data <= jump_crouch_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(7 downto 4);
        --         B_data <= jump_crouch_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(3 downto 0);
        --     when "100" => -- idle1 L
        --         R_data <= idle_1_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(11 downto 8);
        --         G_data <= idle_1_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(7 downto 4);
        --         B_data <= idle_1_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(3 downto 0);
        --     when "101" => -- running1 L
        --         R_data <= running_1_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(11 downto 8);
        --         G_data <= running_1_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(7 downto 4);
        --         B_data <= running_1_L(int_vcount - (int_boundy + 0))(int_hcount - (int_boundx + 0))(3 downto 0);
        --     when others => -- fallback for error handling and checking
        -- R_data <= "0000";
        -- G_data <= "0000";
        -- B_data <= "0000";
        -- end case;
    end process;

end behavioural;