../../VGA/VGA_Vsync_gen_cfg.vhd