../../attack/toplevelattack-structural-cfg.vhd