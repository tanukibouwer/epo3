../../input/input_period_counter_behavioural_cfg.vhd