../../input/input_jump_behavioural_cfg.vhd