../../input/input_toplevel.vhd