../../VGA/VGA_char_animation_fsm_cfg.vhd