configuration p_knockback_calculator_behaviour_cfg of p_knockback_calculator is
   for behaviour
   end for;
end p_knockback_calculator_behaviour_cfg;
