configuration velocity_interpolator_behaviour_cfg of velocity_interpolator is
   for behaviour
   end for;
end velocity_interpolator_behaviour_cfg;
