configuration p_mux_cfg of p_mux is
    for behavioural
    end for;
end configuration p_mux_cfg;