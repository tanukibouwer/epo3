configuration game_state_fsm_cfg of game_state_fsm is
    for behaviour
    end for;
end configuration game_state_fsm_cfg;