../../physics/velocity_interpolator.vhd