../../VGA/VGA_newer_coloring.vhd