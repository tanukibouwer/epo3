../../input/input_driver_behavioural_cfg.vhd