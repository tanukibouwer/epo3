../../memory/m_resethandler.vhd