configuration t_8bregs_rtl_cfg of t_8bregs is
   for rtl
   end for;
end t_8bregs_rtl_cfg;
