../../physics/knockback_calculator.vhd