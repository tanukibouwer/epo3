../../VGA/VGA_char_offset_adder.vhd