../../VGA/VGA_coloring.vhd