
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture routed of chip_toplevel is

  component orientation
    port(clk     : in  std_logic;
         res     : in  std_logic;
         input1  : in  std_logic_vector(7 downto 0);
         input2  : in  std_logic_vector(7 downto 0);
         output1 : out std_logic;
         output2 : out std_logic);
  end component;

  component input_period_counter
    port(clk       : in  std_logic;
         reset     : in  std_logic;
         count_out : out std_logic_vector(3 downto 0));
  end component;

  component DEL01BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL1BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL02BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD1P5BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD12BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD8BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component INVD2BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component IAO21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OR4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component IND3D1BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AO32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component DFKCNQD1BWP7T
    port(CN, CP, D : in std_logic; Q : out std_logic);
  end component;

  component DFQD1BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component EDFKCNQD1BWP7T
    port(CN, CP, D, E : in std_logic; Q : out std_logic);
  end component;

  component AO221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AO211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OA21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component OAI221D1BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component OA211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI33D1BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component AOI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AOI211XD0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OR3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component MAOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AO21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component MAOI222D1BWP7T
    port(A, B, C : in std_logic; ZN : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component INR3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component CKXOR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component FA1D0BWP7T
    port(A, B, CI : in std_logic; CO, S : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component OAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component OAI31D1BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component HA1D0BWP7T
    port(A, B : in std_logic; CO, S : out std_logic);
  end component;

  component AOI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component CKND1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component AOI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component AN4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component CKMUX2D1BWP7T
    port(I0, I1, S : in std_logic; Z : out std_logic);
  end component;

  component IOA21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component XNR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D1P5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component ND4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component IINR4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OA22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component DFD1BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component AO31D1BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component CKND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component XOR3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component OA32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component AOI221D1BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AN3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component AN3D0BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component INR4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component OA221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component IOA21D1BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OA222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; Z : out std_logic);
  end component;

  component OAI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OA33D0BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; Z : out std_logic);
  end component;

  component IND3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component CKAN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component XOR4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component AO32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component AO222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; Z : out std_logic);
  end component;

  component AOI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCND1BWP7T
    port(CN, CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component INVD5BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component DFQD0BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component CKAN2D8BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OA31D1BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component EDFKCND1BWP7T
    port(CN, CP, D, E : in std_logic; Q, QN : out std_logic);
  end component;

  component DFKSND1BWP7T
    port(CP, D, SN : in std_logic; Q, QN : out std_logic);
  end component;

  component AN4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component DFD0BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component CKND10BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component AOI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OAI33D1BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component IND2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component ND3D1BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component OR4XD1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component AOI21D1BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component IIND4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component DFXD1BWP7T
    port(CP, DA, DB, SA : in std_logic; Q, QN : out std_logic);
  end component;

  component IND4D1BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  signal FE_PHN177_char1posyin_1, FE_PHN176_char2velx_9, FE_PHN175_char2vely_3, FE_PHN174_vcountintern_8, FE_PHN173_TL04_driver_pulse_count_0 : std_logic;
  signal FE_PHN172_TL01_CLR1_n_1491, FE_PHN171_TL01_CLR1_char2_sprite_frame_control_frame_count_2, FE_PHN170_TL04_n_15, FE_PHN169_TL01_CLR1_char2_sprite_frame_control_cnt_reset, FE_PHN168_char2posy_7 : std_logic;
  signal FE_PHN167_char1posxin_5, FE_PHN166_TL01_CLR1_char1_sprite_frame_control_cnt_reset, FE_PHN165_char2posx_1, FE_PHN164_char2posx_0, FE_PHN163_TL01_CLR1_char2_sprite_frame_control_frame_count_4 : std_logic;
  signal FE_PHN162_char1posxin_6, FE_PHN161_TL01_CLR1_char1_sprite_frame_control_frame_count_0, FE_PHN160_TL01_SCNR1_hcount_reset, FE_PHN159_char1posyin_1, FE_PHN158_TL01_n_0 : std_logic;
  signal FE_PHN157_ATT1_n_34, FE_PHN156_ATT1_n_26, FE_PHN155_TL04_n_15, FE_PHN154_TL01_CLR1_n_33, FE_PHN153_TL01_CLR1_n_41 : std_logic;
  signal FE_PHN152_TL01_CLR1_n_303, FE_PHN151_TL01_CLR1_n_32, FE_PHN150_TL01_CLR1_n_34, FE_PHN149_TL01_CLR1_n_305, FE_PHN148_ATT1_n_32 : std_logic;
  signal FE_PHN147_TL01_CLR1_n_257, FE_PHN146_ATT1_n_12, FE_PHN145_ATT1_n_35, FE_PHN144_TL01_CLR1_n_733, FE_PHN143_n_73 : std_logic;
  signal FE_PHN142_n_108, FE_PHN141_n_109, FE_PHN140_n_101, FE_PHN139_n_74, FE_PHN138_n_71 : std_logic;
  signal FE_PHN137_n_111, FE_PHN136_n_107, FE_PHN135_n_99, FE_PHN134_n_72, FE_PHN133_n_70 : std_logic;
  signal FE_PHN132_n_75, FE_PHN131_n_105, FE_PHN130_n_98, FE_PHN129_TL04_n_23, FE_PHN128_n_113 : std_logic;
  signal FE_PHN127_n_88, FE_PHN126_ATT1_n_25, FE_PHN125_TL04_n_27, FE_PHN124_char1posx_8, FE_PHN123_char2posx_8 : std_logic;
  signal FE_PHN122_vcountintern_9, FE_PHN121_ATT1_PM2_state2_1, FE_PHN120_ATT1_PM2_state2_0, FE_PHN119_char2posx_6, FE_PHN118_char2perc_1 : std_logic;
  signal FE_PHN117_char2perc_7, FE_PHN116_ATT1_PM2_state1_1, FE_PHN115_ATT1_PM4_state2_1, FE_PHN114_ATT1_PM4_state2_0, FE_PHN113_TL04_driver_state_0 : std_logic;
  signal FE_PHN112_char1perc_7, FE_PHN111_TL01_CLR1_char1_sprite_frame_control_frame_count_2, FE_PHN110_char1perc_0, FE_PHN109_TL01_CLR1_char1_sprite_frame_control_frame_count_3, FE_PHN108_TL01_CLR1_char1_sprite_frame_control_frame_count_0 : std_logic;
  signal FE_PHN107_TL01_CLR1_char2_sprite_frame_control_frame_count_0, FE_PHN106_TL01_CLR1_char1_sprite_frame_control_state_0, FE_PHN105_TL01_CLR1_char1_sprite_frame_control_frame_count_4, FE_PHN104_TL04_driver_state_1, FE_PHN103_TL01_CLR1_char1_sprite_frame_control_state_2 : std_logic;
  signal FE_PHN102_char2perc_0, FE_PHN101_char2posy_2, FE_PHN100_char2posx_3, FE_PHN99_TL01_CLR1_char2_sprite_frame_control_state_2, FE_PHN98_inputsp2_5 : std_logic;
  signal FE_PHN97_char2perc_2, FE_PHN96_TL01_n_1, FE_PHN95_char2posy_0, FE_PHN94_char2posx_1, FE_PHN93_char2posy_6 : std_logic;
  signal FE_PHN92_char2posx_0, FE_PHN91_char2posy_7, FE_PHN90_char2perc_3, FE_PHN89_TL04_n_0, FE_PHN88_TL01_CLR1_char2_sprite_frame_control_state_0 : std_logic;
  signal FE_PHN87_char2velx_9, FE_PHN86_char2vely_3, FE_PHN85_char2posx_2, FE_PHN84_TL01_CLR1_char2_sprite_frame_control_frame_count_3, FE_PHN83_char2posy_3 : std_logic;
  signal FE_PHN82_char2posx_4, FE_PHN81_char2posy_1, FE_PHN80_TL04_driver_pulse_count_0, FE_PHN79_char2posy_4, FE_PHN78_TL04_n_11 : std_logic;
  signal FE_PHN77_char2velx_1, FE_PHN76_char2velx_3, FE_PHN75_char2velx_4, FE_PHN74_TL04_n_13, FE_PHN73_char2velx_0 : std_logic;
  signal FE_PHN72_char2posy_5, FE_PHN71_char2velx_2, FE_PHN70_char2velx_7, FE_PHN69_char1posxin_5, FE_PHN68_TL01_SCNR1_hcount_reset : std_logic;
  signal FE_PHN67_char1posxin_6, FE_PHN66_char2velx_5, FE_PHN65_TL04_n_10, FE_PHN64_TL04_n_12, FE_PHN63_char1posyin_1 : std_logic;
  signal FE_PHN62_TL01_n_0, FE_PHN61_char1velxin_8, FE_PHN60_TL01_CLR1_char2_sprite_frame_control_cnt_reset, FE_PHN59_TL01_CLR1_char1_sprite_frame_control_cnt_reset, FE_PHN58_TL00_WL00_state_1 : std_logic;
  signal FE_PHN57_char1posxin_7, FE_PHN56_char1posxin_2, FE_PHN55_char1posxin_1, FE_PHN54_char1posxin_3, FE_PHN53_TL01_CLR1_n_1 : std_logic;
  signal FE_PHN52_char1posxin_8, FE_PHN51_TL01_CLR1_n_0, FE_PHN50_char1posxin_4, FE_PHN49_char1posxin_0, FE_PHN48_ATT1_n_5 : std_logic;
  signal FE_PHN47_char1posyin_2, FE_PHN46_char1posyin_7, FE_PHN45_char1posyin_6, FE_PHN44_char1posyin_3, FE_PHN43_char1posyin_5 : std_logic;
  signal FE_PHN42_char1posyin_4, FE_PHN41_char1posyin_0, FE_PHN40_char1velyin_9, FE_PHN39_char1velyin_6, FE_PHN38_char1velyin_8 : std_logic;
  signal FE_PHN37_char1velyin_7, FE_PHN36_char1velxin_6, FE_PHN35_char1velyin_1, FE_PHN34_TL01_n_2, FE_PHN33_char1velyin_0 : std_logic;
  signal FE_PHN32_char1velxin_0, FE_PHN31_char1velyin_4, FE_PHN30_char1velyin_2, FE_PHN29_char1velxin_1, FE_PHN28_char1velyin_5 : std_logic;
  signal FE_PHN27_char1velxin_5, FE_PHN26_char1velxin_3, FE_PHN25_char1velxin_2, FE_PHN24_char1velyin_3, FE_PHN23_char1velxin_7 : std_logic;
  signal FE_PHN22_char1velxin_4, FE_PHN21_char1velxin_9, FE_PHN20_TL01_CLR1_char2_sprite_frame_control_new_state_0, FE_PHN19_TL01_CLR1_char1_sprite_frame_control_new_state_0, FE_PHN18_TL01_CLR1_char2_sprite_frame_control_new_state_1 : std_logic;
  signal FE_PHN17_TL01_CLR1_char2_sprite_frame_control_new_state_2, FE_PHN16_TL01_CLR1_char1_sprite_frame_control_new_state_1, FE_PHN15_TL01_CLR1_char1_sprite_frame_control_new_state_2, FE_OFN4_TL00_writeint, FE_OFN3_reset : std_logic;
  signal FE_OFN2_ATT1_n_301, FE_OFN1_TL02_PHS0_sel_0, FE_OFN0_n_6, CTS_18, CTS_17 : std_logic;
  signal CTS_16, CTS_15, FE_DBTN14_reset, FE_DBTN13_char1perc_5, FE_DBTN12_char1perc_4 : std_logic;
  signal FE_DBTN11_char1perc_3, FE_DBTN10_char1perc_1, FE_DBTN9_char2perc_5, FE_DBTN8_char2perc_4, FE_DBTN7_char2perc_3 : std_logic;
  signal FE_DBTN6_char2perc_2, FE_DBTN5_char2perc_1, FE_DBTN4_char2perc_0, FE_DBTN3_char1posx_4, FE_DBTN2_char1posy_3 : std_logic;
  signal FE_DBTN1_char2posx_1, FE_DBTN0_char2posx_0 : std_logic;
  signal dirx2new2 : std_logic_vector(7 downto 0);
  signal dirx1new2 : std_logic_vector(7 downto 0);
  signal char1perctemp : std_logic_vector(7 downto 0);
  signal char2perctemp : std_logic_vector(7 downto 0);
  signal diry1new2 : std_logic_vector(7 downto 0);
  signal diry2new2 : std_logic_vector(7 downto 0);
  signal vcountintern : std_logic_vector(9 downto 0);
  signal diry1new1 : std_logic_vector(7 downto 0);
  signal dirx1new1 : std_logic_vector(7 downto 0);
  signal dirx2new1 : std_logic_vector(7 downto 0);
  signal diry2new1 : std_logic_vector(7 downto 0);
  signal char1perc : std_logic_vector(7 downto 0);
  signal char2perc : std_logic_vector(7 downto 0);
  signal char1posx : std_logic_vector(8 downto 0);
  signal char1posy : std_logic_vector(8 downto 0);
  signal char2posx : std_logic_vector(8 downto 0);
  signal char2posy : std_logic_vector(8 downto 0);
  signal char1velxin : std_logic_vector(9 downto 0);
  signal char1velx : std_logic_vector(9 downto 0);
  signal char1velyin : std_logic_vector(9 downto 0);
  signal char1vely : std_logic_vector(9 downto 0);
  signal char2velx : std_logic_vector(9 downto 0);
  signal char2vely : std_logic_vector(9 downto 0);
  signal char1posxin : std_logic_vector(8 downto 0);
  signal char1posyin : std_logic_vector(8 downto 0);
  signal inputsp1 : std_logic_vector(7 downto 0);
  signal inputsp2 : std_logic_vector(7 downto 0);
  signal char1percin : std_logic_vector(7 downto 0);
  signal char2percin : std_logic_vector(7 downto 0);
  signal hcountintern : std_logic_vector(9 downto 0);
  signal TL04_count : std_logic_vector(3 downto 0);
  signal TL04_deserializer_out_p1 : std_logic_vector(7 downto 0);
  signal TL04_deserializer_out_p2 : std_logic_vector(7 downto 0);
  signal TL01_hcount_int : std_logic_vector(9 downto 0);
  signal ATT1_PM2_state1_0, ATT1_PM2_state1_1, ATT1_PM2_state2_0, ATT1_PM2_state2_1, ATT1_PM3_state1_0 : std_logic;
  signal ATT1_PM3_state1_1, ATT1_PM3_state2_0, ATT1_PM3_state2_1, ATT1_PM4_state1_0, ATT1_PM4_state1_1 : std_logic;
  signal ATT1_PM4_state2_0, ATT1_PM4_state2_1, ATT1_at1a, ATT1_at1b, ATT1_at2a : std_logic;
  signal ATT1_at2b, ATT1_n_0, ATT1_n_1, ATT1_n_3, ATT1_n_4 : std_logic;
  signal ATT1_n_5, ATT1_n_6, ATT1_n_7, ATT1_n_8, ATT1_n_9 : std_logic;
  signal ATT1_n_10, ATT1_n_11, ATT1_n_12, ATT1_n_13, ATT1_n_14 : std_logic;
  signal ATT1_n_15, ATT1_n_16, ATT1_n_17, ATT1_n_18, ATT1_n_19 : std_logic;
  signal ATT1_n_20, ATT1_n_21, ATT1_n_22, ATT1_n_23, ATT1_n_24 : std_logic;
  signal ATT1_n_25, ATT1_n_26, ATT1_n_27, ATT1_n_28, ATT1_n_29 : std_logic;
  signal ATT1_n_30, ATT1_n_31, ATT1_n_32, ATT1_n_33, ATT1_n_34 : std_logic;
  signal ATT1_n_35, ATT1_n_36, ATT1_n_37, ATT1_n_38, ATT1_n_39 : std_logic;
  signal ATT1_n_40, ATT1_n_41, ATT1_n_42, ATT1_n_43, ATT1_n_44 : std_logic;
  signal ATT1_n_47, ATT1_n_49, ATT1_n_50, ATT1_n_51, ATT1_n_53 : std_logic;
  signal ATT1_n_58, ATT1_n_62, ATT1_n_65, ATT1_n_66, ATT1_n_67 : std_logic;
  signal ATT1_n_68, ATT1_n_70, ATT1_n_71, ATT1_n_72, ATT1_n_73 : std_logic;
  signal ATT1_n_74, ATT1_n_75, ATT1_n_76, ATT1_n_77, ATT1_n_78 : std_logic;
  signal ATT1_n_79, ATT1_n_80, ATT1_n_81, ATT1_n_82, ATT1_n_83 : std_logic;
  signal ATT1_n_84, ATT1_n_85, ATT1_n_86, ATT1_n_87, ATT1_n_88 : std_logic;
  signal ATT1_n_89, ATT1_n_90, ATT1_n_91, ATT1_n_92, ATT1_n_93 : std_logic;
  signal ATT1_n_94, ATT1_n_95, ATT1_n_96, ATT1_n_97, ATT1_n_98 : std_logic;
  signal ATT1_n_99, ATT1_n_100, ATT1_n_101, ATT1_n_102, ATT1_n_103 : std_logic;
  signal ATT1_n_104, ATT1_n_105, ATT1_n_106, ATT1_n_107, ATT1_n_108 : std_logic;
  signal ATT1_n_109, ATT1_n_110, ATT1_n_111, ATT1_n_112, ATT1_n_113 : std_logic;
  signal ATT1_n_114, ATT1_n_115, ATT1_n_116, ATT1_n_117, ATT1_n_118 : std_logic;
  signal ATT1_n_119, ATT1_n_120, ATT1_n_121, ATT1_n_122, ATT1_n_123 : std_logic;
  signal ATT1_n_124, ATT1_n_125, ATT1_n_126, ATT1_n_127, ATT1_n_128 : std_logic;
  signal ATT1_n_129, ATT1_n_130, ATT1_n_131, ATT1_n_132, ATT1_n_133 : std_logic;
  signal ATT1_n_134, ATT1_n_135, ATT1_n_136, ATT1_n_137, ATT1_n_138 : std_logic;
  signal ATT1_n_139, ATT1_n_140, ATT1_n_141, ATT1_n_142, ATT1_n_143 : std_logic;
  signal ATT1_n_144, ATT1_n_145, ATT1_n_146, ATT1_n_147, ATT1_n_148 : std_logic;
  signal ATT1_n_149, ATT1_n_150, ATT1_n_151, ATT1_n_152, ATT1_n_153 : std_logic;
  signal ATT1_n_154, ATT1_n_155, ATT1_n_156, ATT1_n_157, ATT1_n_158 : std_logic;
  signal ATT1_n_159, ATT1_n_160, ATT1_n_161, ATT1_n_162, ATT1_n_163 : std_logic;
  signal ATT1_n_164, ATT1_n_165, ATT1_n_166, ATT1_n_167, ATT1_n_168 : std_logic;
  signal ATT1_n_169, ATT1_n_170, ATT1_n_171, ATT1_n_172, ATT1_n_173 : std_logic;
  signal ATT1_n_174, ATT1_n_175, ATT1_n_176, ATT1_n_177, ATT1_n_178 : std_logic;
  signal ATT1_n_179, ATT1_n_180, ATT1_n_181, ATT1_n_182, ATT1_n_183 : std_logic;
  signal ATT1_n_184, ATT1_n_185, ATT1_n_186, ATT1_n_187, ATT1_n_188 : std_logic;
  signal ATT1_n_189, ATT1_n_190, ATT1_n_191, ATT1_n_192, ATT1_n_193 : std_logic;
  signal ATT1_n_194, ATT1_n_195, ATT1_n_196, ATT1_n_197, ATT1_n_198 : std_logic;
  signal ATT1_n_199, ATT1_n_200, ATT1_n_201, ATT1_n_202, ATT1_n_203 : std_logic;
  signal ATT1_n_204, ATT1_n_205, ATT1_n_206, ATT1_n_207, ATT1_n_208 : std_logic;
  signal ATT1_n_209, ATT1_n_210, ATT1_n_211, ATT1_n_212, ATT1_n_213 : std_logic;
  signal ATT1_n_214, ATT1_n_215, ATT1_n_216, ATT1_n_217, ATT1_n_218 : std_logic;
  signal ATT1_n_219, ATT1_n_220, ATT1_n_221, ATT1_n_222, ATT1_n_223 : std_logic;
  signal ATT1_n_224, ATT1_n_225, ATT1_n_226, ATT1_n_227, ATT1_n_228 : std_logic;
  signal ATT1_n_229, ATT1_n_230, ATT1_n_231, ATT1_n_232, ATT1_n_233 : std_logic;
  signal ATT1_n_234, ATT1_n_235, ATT1_n_236, ATT1_n_237, ATT1_n_238 : std_logic;
  signal ATT1_n_239, ATT1_n_240, ATT1_n_241, ATT1_n_242, ATT1_n_243 : std_logic;
  signal ATT1_n_244, ATT1_n_245, ATT1_n_246, ATT1_n_247, ATT1_n_248 : std_logic;
  signal ATT1_n_249, ATT1_n_250, ATT1_n_251, ATT1_n_252, ATT1_n_253 : std_logic;
  signal ATT1_n_254, ATT1_n_255, ATT1_n_256, ATT1_n_257, ATT1_n_258 : std_logic;
  signal ATT1_n_259, ATT1_n_260, ATT1_n_261, ATT1_n_262, ATT1_n_263 : std_logic;
  signal ATT1_n_264, ATT1_n_265, ATT1_n_266, ATT1_n_267, ATT1_n_268 : std_logic;
  signal ATT1_n_269, ATT1_n_270, ATT1_n_271, ATT1_n_272, ATT1_n_273 : std_logic;
  signal ATT1_n_274, ATT1_n_275, ATT1_n_276, ATT1_n_277, ATT1_n_278 : std_logic;
  signal ATT1_n_279, ATT1_n_280, ATT1_n_281, ATT1_n_282, ATT1_n_283 : std_logic;
  signal ATT1_n_284, ATT1_n_285, ATT1_n_286, ATT1_n_287, ATT1_n_288 : std_logic;
  signal ATT1_n_289, ATT1_n_290, ATT1_n_291, ATT1_n_292, ATT1_n_293 : std_logic;
  signal ATT1_n_294, ATT1_n_295, ATT1_n_296, ATT1_n_297, ATT1_n_298 : std_logic;
  signal ATT1_n_299, ATT1_n_300, ATT1_n_301, ATT1_n_302, ATT1_n_303 : std_logic;
  signal ATT1_n_304, ATT1_n_305, ATT1_n_306, ATT1_n_307, ATT1_n_308 : std_logic;
  signal ATT1_n_309, ATT1_n_310, ATT1_n_311, ATT1_n_312, ATT1_n_313 : std_logic;
  signal ATT1_n_314, ATT1_n_315, ATT1_n_316, ATT1_n_317, ATT1_n_318 : std_logic;
  signal ATT1_n_319, ATT1_n_320, ATT1_n_321, ATT1_n_322, ATT1_n_323 : std_logic;
  signal ATT1_n_324, ATT1_n_325, ATT1_n_326, ATT1_n_327, ATT1_n_328 : std_logic;
  signal ATT1_n_329, ATT1_n_330, ATT1_n_331, ATT1_n_332, ATT1_n_333 : std_logic;
  signal ATT1_n_334, ATT1_n_335, ATT1_n_336, ATT1_n_337, ATT1_n_338 : std_logic;
  signal ATT1_n_339, ATT1_n_340, ATT1_n_341, ATT1_n_342, ATT1_n_343 : std_logic;
  signal ATT1_n_344, ATT1_n_345, ATT1_n_346, ATT1_n_347, ATT1_n_348 : std_logic;
  signal ATT1_n_349, ATT1_n_350, ATT1_n_351, ATT1_n_352, ATT1_n_353 : std_logic;
  signal ATT1_n_354, ATT1_n_355, ATT1_n_356, ATT1_n_357, ATT1_n_358 : std_logic;
  signal ATT1_n_359, ATT1_n_360, ATT1_n_361, ATT1_n_362, ATT1_n_363 : std_logic;
  signal ATT1_n_364, ATT1_n_365, ATT1_n_366, ATT1_n_367, ATT1_n_368 : std_logic;
  signal ATT1_n_369, ATT1_n_370, ATT1_n_371, ATT1_n_372, ATT1_n_373 : std_logic;
  signal ATT1_n_374, ATT1_n_375, ATT1_n_376, ATT1_n_377, ATT1_n_378 : std_logic;
  signal ATT1_n_379, ATT1_n_380, ATT1_n_381, ATT1_n_382, ATT1_n_383 : std_logic;
  signal ATT1_n_384, ATT1_n_385, ATT1_n_386, ATT1_n_387, ATT1_n_388 : std_logic;
  signal ATT1_n_389, ATT1_n_390, ATT1_n_391, ATT1_n_392, ATT1_n_393 : std_logic;
  signal ATT1_n_394, ATT1_n_395, ATT1_n_396, ATT1_n_397, ATT1_n_398 : std_logic;
  signal ATT1_n_399, ATT1_n_400, ATT1_n_401, ATT1_n_402, ATT1_n_403 : std_logic;
  signal ATT1_n_404, ATT1_n_405, ATT1_n_406, ATT1_n_407, ATT1_n_408 : std_logic;
  signal ATT1_n_409, ATT1_n_410, ATT1_n_411, ATT1_n_412, ATT1_n_413 : std_logic;
  signal ATT1_n_414, ATT1_n_415, ATT1_n_416, ATT1_n_417, ATT1_n_418 : std_logic;
  signal ATT1_n_419, ATT1_n_420, ATT1_n_421, ATT1_n_422, ATT1_n_423 : std_logic;
  signal ATT1_n_424, ATT1_n_425, ATT1_n_426, ATT1_n_427, ATT1_n_428 : std_logic;
  signal ATT1_n_429, ATT1_n_430, ATT1_n_431, ATT1_n_432, ATT1_n_433 : std_logic;
  signal ATT1_n_434, ATT1_n_435, ATT1_n_436, ATT1_n_437, ATT1_n_438 : std_logic;
  signal ATT1_n_439, ATT1_n_440, ATT1_n_441, ATT1_n_442, ATT1_n_443 : std_logic;
  signal ATT1_n_444, ATT1_n_445, ATT1_n_446, ATT1_n_447, ATT1_n_448 : std_logic;
  signal ATT1_n_449, ATT1_n_450, ATT1_n_451, ATT1_n_452, ATT1_n_453 : std_logic;
  signal ATT1_n_454, ATT1_n_455, ATT1_n_456, ATT1_n_457, ATT1_n_458 : std_logic;
  signal ATT1_n_459, ATT1_n_460, ATT1_n_461, ATT1_n_462, ATT1_n_463 : std_logic;
  signal ATT1_n_464, ATT1_n_465, ATT1_n_466, ATT1_n_467, ATT1_n_468 : std_logic;
  signal ATT1_n_469, ATT1_n_470, ATT1_n_471, ATT1_n_472, ATT1_n_473 : std_logic;
  signal ATT1_n_474, ATT1_n_475, ATT1_n_476, ATT1_n_477, ATT1_n_478 : std_logic;
  signal ATT1_n_479, ATT1_n_480, ATT1_n_481, ATT1_n_482, ATT1_n_483 : std_logic;
  signal ATT1_n_484, ATT1_n_485, ATT1_n_486, ATT1_n_487, ATT1_n_488 : std_logic;
  signal ATT1_n_489, ATT1_n_490, ATT1_n_491, ATT1_n_492, ATT1_n_493 : std_logic;
  signal ATT1_n_494, ATT1_n_495, ATT1_n_496, ATT1_n_497, ATT1_n_498 : std_logic;
  signal ATT1_n_499, ATT1_n_500, ATT1_n_501, ATT1_n_502, ATT1_n_503 : std_logic;
  signal ATT1_n_504, ATT1_n_505, ATT1_n_506, ATT1_n_507, ATT1_n_508 : std_logic;
  signal ATT1_n_509, ATT1_n_510, ATT1_n_511, ATT1_n_512, ATT1_n_513 : std_logic;
  signal ATT1_n_514, ATT1_n_515, ATT1_n_516, ATT1_n_517, ATT1_n_518 : std_logic;
  signal ATT1_n_519, ATT1_n_520, ATT1_n_521, ATT1_n_522, ATT1_n_523 : std_logic;
  signal ATT1_n_524, ATT1_n_525, ATT1_n_526, ATT1_n_527, ATT1_n_528 : std_logic;
  signal ATT1_n_529, ATT1_n_530, ATT1_n_531, ATT1_n_532, ATT1_n_533 : std_logic;
  signal ATT1_n_534, ATT1_n_535, ATT1_n_536, ATT1_n_537, ATT1_n_538 : std_logic;
  signal ATT1_n_539, ATT1_n_540, ATT1_n_541, ATT1_n_542, ATT1_n_543 : std_logic;
  signal ATT1_n_544, ATT1_n_545, ATT1_n_546, ATT1_n_547, ATT1_n_548 : std_logic;
  signal ATT1_n_549, ATT1_n_550, ATT1_n_551, ATT1_n_552, ATT1_n_553 : std_logic;
  signal ATT1_n_554, ATT1_n_555, ATT1_n_556, ATT1_n_557, ATT1_n_558 : std_logic;
  signal ATT1_n_559, ATT1_n_560, ATT1_n_561, ATT1_n_562, ATT1_n_563 : std_logic;
  signal ATT1_n_564, ATT1_n_565, ATT1_n_566, ATT1_n_567, ATT1_n_568 : std_logic;
  signal ATT1_n_569, ATT1_n_570, ATT1_n_571, ATT1_n_572, ATT1_n_573 : std_logic;
  signal ATT1_n_574, ATT1_n_575, ATT1_n_576, ATT1_n_577, ATT1_n_578 : std_logic;
  signal ATT1_n_579, ATT1_n_580, ATT1_n_581, ATT1_n_582, ATT1_n_583 : std_logic;
  signal ATT1_n_584, ATT1_n_585, ATT1_n_586, ATT1_n_587, ATT1_n_588 : std_logic;
  signal ATT1_n_589, ATT1_n_590, ATT1_n_591, ATT1_n_592, ATT1_n_593 : std_logic;
  signal ATT1_n_594, ATT1_n_595, ATT1_n_596, ATT1_n_597, ATT1_n_598 : std_logic;
  signal ATT1_n_599, ATT1_n_600, ATT1_n_601, ATT1_n_602, ATT1_n_603 : std_logic;
  signal ATT1_n_604, ATT1_n_605, ATT1_n_606, ATT1_n_607, ATT1_n_608 : std_logic;
  signal ATT1_n_609, ATT1_n_610, ATT1_n_611, ATT1_n_612, ATT1_n_613 : std_logic;
  signal ATT1_n_614, ATT1_n_615, ATT1_n_616, ATT1_n_617, ATT1_n_618 : std_logic;
  signal ATT1_n_619, ATT1_n_620, ATT1_n_621, ATT1_n_622, ATT1_n_623 : std_logic;
  signal ATT1_n_624, ATT1_n_625, ATT1_n_626, ATT1_n_627, ATT1_n_628 : std_logic;
  signal ATT1_n_629, ATT1_n_630, ATT1_n_631, ATT1_n_632, ATT1_n_633 : std_logic;
  signal ATT1_n_634, ATT1_n_635, ATT1_n_636, ATT1_n_637, ATT1_n_638 : std_logic;
  signal ATT1_n_639, ATT1_n_640, ATT1_n_641, ATT1_n_642, ATT1_n_643 : std_logic;
  signal ATT1_n_644, ATT1_n_645, ATT1_n_646, ATT1_n_647, ATT1_n_648 : std_logic;
  signal ATT1_n_649, ATT1_n_650, ATT1_n_651, ATT1_n_652, ATT1_n_653 : std_logic;
  signal ATT1_n_654, ATT1_n_655, ATT1_n_656, ATT1_n_657, ATT1_n_658 : std_logic;
  signal ATT1_n_659, ATT1_n_660, ATT1_n_661, ATT1_n_662, ATT1_n_663 : std_logic;
  signal ATT1_n_664, ATT1_n_665, ATT1_n_666, ATT1_n_667, ATT1_n_668 : std_logic;
  signal ATT1_n_669, ATT1_n_670, ATT1_n_671, ATT1_n_672, ATT1_n_673 : std_logic;
  signal ATT1_n_674, ATT1_n_675, ATT1_n_676, ATT1_n_677, ATT1_n_678 : std_logic;
  signal ATT1_n_679, ATT1_n_680, ATT1_n_681, ATT1_n_682, ATT1_n_683 : std_logic;
  signal ATT1_n_684, ATT1_n_685, ATT1_n_686, ATT1_n_687, ATT1_n_688 : std_logic;
  signal ATT1_n_689, ATT1_n_690, ATT1_n_691, ATT1_n_692, ATT1_n_693 : std_logic;
  signal ATT1_n_694, ATT1_n_695, ATT1_n_696, ATT1_n_697, ATT1_n_698 : std_logic;
  signal ATT1_n_699, ATT1_n_700, ATT1_n_701, ATT1_n_702, ATT1_n_703 : std_logic;
  signal ATT1_n_704, ATT1_n_705, ATT1_n_706, ATT1_n_707, ATT1_n_708 : std_logic;
  signal ATT1_n_709, ATT1_n_710, ATT1_n_711, ATT1_n_712, ATT1_n_713 : std_logic;
  signal ATT1_n_714, ATT1_n_715, ATT1_n_716, ATT1_n_717, ATT1_n_718 : std_logic;
  signal ATT1_n_719, ATT1_n_720, ATT1_n_721, ATT1_n_722, ATT1_n_723 : std_logic;
  signal ATT1_n_724, ATT1_n_725, ATT1_n_726, ATT1_n_727, ATT1_n_728 : std_logic;
  signal ATT1_n_729, ATT1_n_730, ATT1_n_731, ATT1_n_732, ATT1_n_733 : std_logic;
  signal ATT1_n_734, ATT1_n_735, ATT1_n_736, ATT1_n_737, ATT1_n_738 : std_logic;
  signal ATT1_n_739, ATT1_n_740, ATT1_n_741, ATT1_n_742, ATT1_n_743 : std_logic;
  signal ATT1_n_744, ATT1_n_745, ATT1_n_746, ATT1_n_747, ATT1_n_748 : std_logic;
  signal ATT1_n_749, ATT1_n_750, ATT1_n_751, ATT1_n_752, ATT1_n_753 : std_logic;
  signal ATT1_n_754, ATT1_n_755, ATT1_n_756, ATT1_n_757, ATT1_n_758 : std_logic;
  signal ATT1_n_759, ATT1_n_817, ATT1_n_818, ATT1_n_827, ATT1_n_828 : std_logic;
  signal TL00_WL00_state_1, TL00_writeint, TL01_CLR1_char1_sprite_frame_control_cnt_reset, TL01_CLR1_char1_sprite_frame_control_frame_count_0, TL01_CLR1_char1_sprite_frame_control_frame_count_1 : std_logic;
  signal TL01_CLR1_char1_sprite_frame_control_frame_count_2, TL01_CLR1_char1_sprite_frame_control_frame_count_3, TL01_CLR1_char1_sprite_frame_control_frame_count_4, TL01_CLR1_char1_sprite_frame_control_new_state_0, TL01_CLR1_char1_sprite_frame_control_new_state_1 : std_logic;
  signal TL01_CLR1_char1_sprite_frame_control_new_state_2, TL01_CLR1_char1_sprite_frame_control_state_0, TL01_CLR1_char1_sprite_frame_control_state_1, TL01_CLR1_char1_sprite_frame_control_state_2, TL01_CLR1_char1_sprite_sprite_0 : std_logic;
  signal TL01_CLR1_char1_sprite_sprite_1, TL01_CLR1_char2_sprite_frame_control_cnt_reset, TL01_CLR1_char2_sprite_frame_control_frame_count_0, TL01_CLR1_char2_sprite_frame_control_frame_count_1, TL01_CLR1_char2_sprite_frame_control_frame_count_2 : std_logic;
  signal TL01_CLR1_char2_sprite_frame_control_frame_count_3, TL01_CLR1_char2_sprite_frame_control_frame_count_4, TL01_CLR1_char2_sprite_frame_control_new_state_0, TL01_CLR1_char2_sprite_frame_control_new_state_1, TL01_CLR1_char2_sprite_frame_control_new_state_2 : std_logic;
  signal TL01_CLR1_char2_sprite_frame_control_state_0, TL01_CLR1_char2_sprite_frame_control_state_1, TL01_CLR1_char2_sprite_frame_control_state_2, TL01_CLR1_char2_sprite_sprite_0, TL01_CLR1_char2_sprite_sprite_1 : std_logic;
  signal TL01_CLR1_n_0, TL01_CLR1_n_1, TL01_CLR1_n_2, TL01_CLR1_n_3, TL01_CLR1_n_5 : std_logic;
  signal TL01_CLR1_n_6, TL01_CLR1_n_9, TL01_CLR1_n_10, TL01_CLR1_n_11, TL01_CLR1_n_12 : std_logic;
  signal TL01_CLR1_n_13, TL01_CLR1_n_14, TL01_CLR1_n_15, TL01_CLR1_n_16, TL01_CLR1_n_17 : std_logic;
  signal TL01_CLR1_n_18, TL01_CLR1_n_19, TL01_CLR1_n_20, TL01_CLR1_n_21, TL01_CLR1_n_22 : std_logic;
  signal TL01_CLR1_n_23, TL01_CLR1_n_24, TL01_CLR1_n_25, TL01_CLR1_n_26, TL01_CLR1_n_27 : std_logic;
  signal TL01_CLR1_n_28, TL01_CLR1_n_29, TL01_CLR1_n_30, TL01_CLR1_n_31, TL01_CLR1_n_32 : std_logic;
  signal TL01_CLR1_n_33, TL01_CLR1_n_34, TL01_CLR1_n_35, TL01_CLR1_n_36, TL01_CLR1_n_37 : std_logic;
  signal TL01_CLR1_n_38, TL01_CLR1_n_39, TL01_CLR1_n_40, TL01_CLR1_n_41, TL01_CLR1_n_42 : std_logic;
  signal TL01_CLR1_n_43, TL01_CLR1_n_44, TL01_CLR1_n_45, TL01_CLR1_n_46, TL01_CLR1_n_47 : std_logic;
  signal TL01_CLR1_n_48, TL01_CLR1_n_49, TL01_CLR1_n_50, TL01_CLR1_n_51, TL01_CLR1_n_52 : std_logic;
  signal TL01_CLR1_n_53, TL01_CLR1_n_54, TL01_CLR1_n_55, TL01_CLR1_n_56, TL01_CLR1_n_57 : std_logic;
  signal TL01_CLR1_n_59, TL01_CLR1_n_60, TL01_CLR1_n_61, TL01_CLR1_n_65, TL01_CLR1_n_66 : std_logic;
  signal TL01_CLR1_n_68, TL01_CLR1_n_69, TL01_CLR1_n_71, TL01_CLR1_n_72, TL01_CLR1_n_73 : std_logic;
  signal TL01_CLR1_n_74, TL01_CLR1_n_75, TL01_CLR1_n_77, TL01_CLR1_n_81, TL01_CLR1_n_82 : std_logic;
  signal TL01_CLR1_n_83, TL01_CLR1_n_84, TL01_CLR1_n_85, TL01_CLR1_n_86, TL01_CLR1_n_87 : std_logic;
  signal TL01_CLR1_n_90, TL01_CLR1_n_92, TL01_CLR1_n_95, TL01_CLR1_n_97, TL01_CLR1_n_98 : std_logic;
  signal TL01_CLR1_n_99, TL01_CLR1_n_100, TL01_CLR1_n_101, TL01_CLR1_n_102, TL01_CLR1_n_103 : std_logic;
  signal TL01_CLR1_n_104, TL01_CLR1_n_105, TL01_CLR1_n_106, TL01_CLR1_n_107, TL01_CLR1_n_108 : std_logic;
  signal TL01_CLR1_n_109, TL01_CLR1_n_110, TL01_CLR1_n_111, TL01_CLR1_n_112, TL01_CLR1_n_113 : std_logic;
  signal TL01_CLR1_n_114, TL01_CLR1_n_115, TL01_CLR1_n_116, TL01_CLR1_n_117, TL01_CLR1_n_118 : std_logic;
  signal TL01_CLR1_n_119, TL01_CLR1_n_120, TL01_CLR1_n_121, TL01_CLR1_n_123, TL01_CLR1_n_124 : std_logic;
  signal TL01_CLR1_n_125, TL01_CLR1_n_126, TL01_CLR1_n_127, TL01_CLR1_n_128, TL01_CLR1_n_129 : std_logic;
  signal TL01_CLR1_n_130, TL01_CLR1_n_131, TL01_CLR1_n_132, TL01_CLR1_n_133, TL01_CLR1_n_134 : std_logic;
  signal TL01_CLR1_n_135, TL01_CLR1_n_136, TL01_CLR1_n_137, TL01_CLR1_n_138, TL01_CLR1_n_139 : std_logic;
  signal TL01_CLR1_n_140, TL01_CLR1_n_141, TL01_CLR1_n_142, TL01_CLR1_n_143, TL01_CLR1_n_144 : std_logic;
  signal TL01_CLR1_n_145, TL01_CLR1_n_146, TL01_CLR1_n_147, TL01_CLR1_n_148, TL01_CLR1_n_149 : std_logic;
  signal TL01_CLR1_n_150, TL01_CLR1_n_151, TL01_CLR1_n_152, TL01_CLR1_n_153, TL01_CLR1_n_154 : std_logic;
  signal TL01_CLR1_n_155, TL01_CLR1_n_156, TL01_CLR1_n_157, TL01_CLR1_n_158, TL01_CLR1_n_159 : std_logic;
  signal TL01_CLR1_n_160, TL01_CLR1_n_161, TL01_CLR1_n_162, TL01_CLR1_n_163, TL01_CLR1_n_164 : std_logic;
  signal TL01_CLR1_n_165, TL01_CLR1_n_166, TL01_CLR1_n_167, TL01_CLR1_n_168, TL01_CLR1_n_169 : std_logic;
  signal TL01_CLR1_n_170, TL01_CLR1_n_171, TL01_CLR1_n_172, TL01_CLR1_n_173, TL01_CLR1_n_174 : std_logic;
  signal TL01_CLR1_n_175, TL01_CLR1_n_176, TL01_CLR1_n_177, TL01_CLR1_n_178, TL01_CLR1_n_179 : std_logic;
  signal TL01_CLR1_n_180, TL01_CLR1_n_181, TL01_CLR1_n_182, TL01_CLR1_n_183, TL01_CLR1_n_184 : std_logic;
  signal TL01_CLR1_n_185, TL01_CLR1_n_186, TL01_CLR1_n_187, TL01_CLR1_n_188, TL01_CLR1_n_189 : std_logic;
  signal TL01_CLR1_n_190, TL01_CLR1_n_191, TL01_CLR1_n_192, TL01_CLR1_n_193, TL01_CLR1_n_194 : std_logic;
  signal TL01_CLR1_n_195, TL01_CLR1_n_196, TL01_CLR1_n_197, TL01_CLR1_n_198, TL01_CLR1_n_199 : std_logic;
  signal TL01_CLR1_n_200, TL01_CLR1_n_201, TL01_CLR1_n_202, TL01_CLR1_n_203, TL01_CLR1_n_204 : std_logic;
  signal TL01_CLR1_n_205, TL01_CLR1_n_206, TL01_CLR1_n_207, TL01_CLR1_n_208, TL01_CLR1_n_209 : std_logic;
  signal TL01_CLR1_n_211, TL01_CLR1_n_212, TL01_CLR1_n_213, TL01_CLR1_n_214, TL01_CLR1_n_215 : std_logic;
  signal TL01_CLR1_n_216, TL01_CLR1_n_217, TL01_CLR1_n_218, TL01_CLR1_n_219, TL01_CLR1_n_220 : std_logic;
  signal TL01_CLR1_n_221, TL01_CLR1_n_222, TL01_CLR1_n_223, TL01_CLR1_n_224, TL01_CLR1_n_225 : std_logic;
  signal TL01_CLR1_n_226, TL01_CLR1_n_227, TL01_CLR1_n_228, TL01_CLR1_n_229, TL01_CLR1_n_230 : std_logic;
  signal TL01_CLR1_n_231, TL01_CLR1_n_232, TL01_CLR1_n_233, TL01_CLR1_n_234, TL01_CLR1_n_235 : std_logic;
  signal TL01_CLR1_n_236, TL01_CLR1_n_237, TL01_CLR1_n_238, TL01_CLR1_n_239, TL01_CLR1_n_240 : std_logic;
  signal TL01_CLR1_n_241, TL01_CLR1_n_242, TL01_CLR1_n_245, TL01_CLR1_n_246, TL01_CLR1_n_247 : std_logic;
  signal TL01_CLR1_n_248, TL01_CLR1_n_249, TL01_CLR1_n_250, TL01_CLR1_n_251, TL01_CLR1_n_252 : std_logic;
  signal TL01_CLR1_n_253, TL01_CLR1_n_254, TL01_CLR1_n_255, TL01_CLR1_n_256, TL01_CLR1_n_257 : std_logic;
  signal TL01_CLR1_n_258, TL01_CLR1_n_259, TL01_CLR1_n_260, TL01_CLR1_n_261, TL01_CLR1_n_262 : std_logic;
  signal TL01_CLR1_n_263, TL01_CLR1_n_264, TL01_CLR1_n_265, TL01_CLR1_n_266, TL01_CLR1_n_267 : std_logic;
  signal TL01_CLR1_n_268, TL01_CLR1_n_269, TL01_CLR1_n_270, TL01_CLR1_n_271, TL01_CLR1_n_272 : std_logic;
  signal TL01_CLR1_n_273, TL01_CLR1_n_274, TL01_CLR1_n_275, TL01_CLR1_n_276, TL01_CLR1_n_277 : std_logic;
  signal TL01_CLR1_n_278, TL01_CLR1_n_279, TL01_CLR1_n_280, TL01_CLR1_n_281, TL01_CLR1_n_282 : std_logic;
  signal TL01_CLR1_n_283, TL01_CLR1_n_284, TL01_CLR1_n_285, TL01_CLR1_n_286, TL01_CLR1_n_287 : std_logic;
  signal TL01_CLR1_n_288, TL01_CLR1_n_289, TL01_CLR1_n_290, TL01_CLR1_n_291, TL01_CLR1_n_292 : std_logic;
  signal TL01_CLR1_n_293, TL01_CLR1_n_294, TL01_CLR1_n_295, TL01_CLR1_n_296, TL01_CLR1_n_297 : std_logic;
  signal TL01_CLR1_n_298, TL01_CLR1_n_299, TL01_CLR1_n_300, TL01_CLR1_n_301, TL01_CLR1_n_302 : std_logic;
  signal TL01_CLR1_n_303, TL01_CLR1_n_304, TL01_CLR1_n_305, TL01_CLR1_n_306, TL01_CLR1_n_307 : std_logic;
  signal TL01_CLR1_n_308, TL01_CLR1_n_309, TL01_CLR1_n_310, TL01_CLR1_n_311, TL01_CLR1_n_312 : std_logic;
  signal TL01_CLR1_n_313, TL01_CLR1_n_314, TL01_CLR1_n_315, TL01_CLR1_n_316, TL01_CLR1_n_317 : std_logic;
  signal TL01_CLR1_n_318, TL01_CLR1_n_319, TL01_CLR1_n_320, TL01_CLR1_n_321, TL01_CLR1_n_322 : std_logic;
  signal TL01_CLR1_n_323, TL01_CLR1_n_324, TL01_CLR1_n_325, TL01_CLR1_n_326, TL01_CLR1_n_327 : std_logic;
  signal TL01_CLR1_n_328, TL01_CLR1_n_329, TL01_CLR1_n_330, TL01_CLR1_n_331, TL01_CLR1_n_332 : std_logic;
  signal TL01_CLR1_n_333, TL01_CLR1_n_334, TL01_CLR1_n_335, TL01_CLR1_n_336, TL01_CLR1_n_337 : std_logic;
  signal TL01_CLR1_n_338, TL01_CLR1_n_339, TL01_CLR1_n_340, TL01_CLR1_n_341, TL01_CLR1_n_342 : std_logic;
  signal TL01_CLR1_n_343, TL01_CLR1_n_345, TL01_CLR1_n_346, TL01_CLR1_n_347, TL01_CLR1_n_348 : std_logic;
  signal TL01_CLR1_n_349, TL01_CLR1_n_350, TL01_CLR1_n_351, TL01_CLR1_n_352, TL01_CLR1_n_353 : std_logic;
  signal TL01_CLR1_n_354, TL01_CLR1_n_355, TL01_CLR1_n_356, TL01_CLR1_n_357, TL01_CLR1_n_358 : std_logic;
  signal TL01_CLR1_n_359, TL01_CLR1_n_360, TL01_CLR1_n_361, TL01_CLR1_n_362, TL01_CLR1_n_363 : std_logic;
  signal TL01_CLR1_n_364, TL01_CLR1_n_365, TL01_CLR1_n_366, TL01_CLR1_n_367, TL01_CLR1_n_368 : std_logic;
  signal TL01_CLR1_n_369, TL01_CLR1_n_370, TL01_CLR1_n_371, TL01_CLR1_n_372, TL01_CLR1_n_373 : std_logic;
  signal TL01_CLR1_n_374, TL01_CLR1_n_375, TL01_CLR1_n_376, TL01_CLR1_n_377, TL01_CLR1_n_378 : std_logic;
  signal TL01_CLR1_n_379, TL01_CLR1_n_380, TL01_CLR1_n_381, TL01_CLR1_n_382, TL01_CLR1_n_383 : std_logic;
  signal TL01_CLR1_n_384, TL01_CLR1_n_385, TL01_CLR1_n_386, TL01_CLR1_n_387, TL01_CLR1_n_388 : std_logic;
  signal TL01_CLR1_n_389, TL01_CLR1_n_390, TL01_CLR1_n_391, TL01_CLR1_n_392, TL01_CLR1_n_393 : std_logic;
  signal TL01_CLR1_n_394, TL01_CLR1_n_395, TL01_CLR1_n_396, TL01_CLR1_n_397, TL01_CLR1_n_398 : std_logic;
  signal TL01_CLR1_n_399, TL01_CLR1_n_400, TL01_CLR1_n_401, TL01_CLR1_n_402, TL01_CLR1_n_403 : std_logic;
  signal TL01_CLR1_n_404, TL01_CLR1_n_405, TL01_CLR1_n_406, TL01_CLR1_n_407, TL01_CLR1_n_408 : std_logic;
  signal TL01_CLR1_n_409, TL01_CLR1_n_410, TL01_CLR1_n_411, TL01_CLR1_n_412, TL01_CLR1_n_413 : std_logic;
  signal TL01_CLR1_n_414, TL01_CLR1_n_415, TL01_CLR1_n_416, TL01_CLR1_n_417, TL01_CLR1_n_418 : std_logic;
  signal TL01_CLR1_n_419, TL01_CLR1_n_420, TL01_CLR1_n_421, TL01_CLR1_n_422, TL01_CLR1_n_423 : std_logic;
  signal TL01_CLR1_n_424, TL01_CLR1_n_425, TL01_CLR1_n_426, TL01_CLR1_n_427, TL01_CLR1_n_428 : std_logic;
  signal TL01_CLR1_n_429, TL01_CLR1_n_430, TL01_CLR1_n_431, TL01_CLR1_n_432, TL01_CLR1_n_433 : std_logic;
  signal TL01_CLR1_n_434, TL01_CLR1_n_435, TL01_CLR1_n_436, TL01_CLR1_n_437, TL01_CLR1_n_438 : std_logic;
  signal TL01_CLR1_n_439, TL01_CLR1_n_440, TL01_CLR1_n_441, TL01_CLR1_n_442, TL01_CLR1_n_443 : std_logic;
  signal TL01_CLR1_n_444, TL01_CLR1_n_445, TL01_CLR1_n_446, TL01_CLR1_n_447, TL01_CLR1_n_448 : std_logic;
  signal TL01_CLR1_n_449, TL01_CLR1_n_450, TL01_CLR1_n_451, TL01_CLR1_n_452, TL01_CLR1_n_453 : std_logic;
  signal TL01_CLR1_n_454, TL01_CLR1_n_455, TL01_CLR1_n_456, TL01_CLR1_n_457, TL01_CLR1_n_458 : std_logic;
  signal TL01_CLR1_n_459, TL01_CLR1_n_460, TL01_CLR1_n_461, TL01_CLR1_n_462, TL01_CLR1_n_463 : std_logic;
  signal TL01_CLR1_n_464, TL01_CLR1_n_465, TL01_CLR1_n_466, TL01_CLR1_n_467, TL01_CLR1_n_468 : std_logic;
  signal TL01_CLR1_n_469, TL01_CLR1_n_470, TL01_CLR1_n_471, TL01_CLR1_n_472, TL01_CLR1_n_473 : std_logic;
  signal TL01_CLR1_n_474, TL01_CLR1_n_475, TL01_CLR1_n_476, TL01_CLR1_n_477, TL01_CLR1_n_478 : std_logic;
  signal TL01_CLR1_n_479, TL01_CLR1_n_480, TL01_CLR1_n_481, TL01_CLR1_n_482, TL01_CLR1_n_483 : std_logic;
  signal TL01_CLR1_n_484, TL01_CLR1_n_485, TL01_CLR1_n_486, TL01_CLR1_n_487, TL01_CLR1_n_488 : std_logic;
  signal TL01_CLR1_n_489, TL01_CLR1_n_490, TL01_CLR1_n_491, TL01_CLR1_n_492, TL01_CLR1_n_493 : std_logic;
  signal TL01_CLR1_n_494, TL01_CLR1_n_495, TL01_CLR1_n_496, TL01_CLR1_n_497, TL01_CLR1_n_498 : std_logic;
  signal TL01_CLR1_n_499, TL01_CLR1_n_500, TL01_CLR1_n_501, TL01_CLR1_n_502, TL01_CLR1_n_503 : std_logic;
  signal TL01_CLR1_n_504, TL01_CLR1_n_505, TL01_CLR1_n_506, TL01_CLR1_n_507, TL01_CLR1_n_508 : std_logic;
  signal TL01_CLR1_n_509, TL01_CLR1_n_510, TL01_CLR1_n_511, TL01_CLR1_n_512, TL01_CLR1_n_513 : std_logic;
  signal TL01_CLR1_n_514, TL01_CLR1_n_515, TL01_CLR1_n_516, TL01_CLR1_n_517, TL01_CLR1_n_518 : std_logic;
  signal TL01_CLR1_n_519, TL01_CLR1_n_520, TL01_CLR1_n_521, TL01_CLR1_n_522, TL01_CLR1_n_523 : std_logic;
  signal TL01_CLR1_n_524, TL01_CLR1_n_525, TL01_CLR1_n_526, TL01_CLR1_n_527, TL01_CLR1_n_528 : std_logic;
  signal TL01_CLR1_n_529, TL01_CLR1_n_530, TL01_CLR1_n_531, TL01_CLR1_n_532, TL01_CLR1_n_533 : std_logic;
  signal TL01_CLR1_n_534, TL01_CLR1_n_535, TL01_CLR1_n_536, TL01_CLR1_n_537, TL01_CLR1_n_538 : std_logic;
  signal TL01_CLR1_n_539, TL01_CLR1_n_540, TL01_CLR1_n_541, TL01_CLR1_n_542, TL01_CLR1_n_543 : std_logic;
  signal TL01_CLR1_n_544, TL01_CLR1_n_545, TL01_CLR1_n_546, TL01_CLR1_n_547, TL01_CLR1_n_548 : std_logic;
  signal TL01_CLR1_n_549, TL01_CLR1_n_550, TL01_CLR1_n_551, TL01_CLR1_n_552, TL01_CLR1_n_553 : std_logic;
  signal TL01_CLR1_n_554, TL01_CLR1_n_555, TL01_CLR1_n_556, TL01_CLR1_n_557, TL01_CLR1_n_558 : std_logic;
  signal TL01_CLR1_n_559, TL01_CLR1_n_560, TL01_CLR1_n_561, TL01_CLR1_n_562, TL01_CLR1_n_563 : std_logic;
  signal TL01_CLR1_n_564, TL01_CLR1_n_565, TL01_CLR1_n_566, TL01_CLR1_n_567, TL01_CLR1_n_568 : std_logic;
  signal TL01_CLR1_n_569, TL01_CLR1_n_570, TL01_CLR1_n_571, TL01_CLR1_n_572, TL01_CLR1_n_573 : std_logic;
  signal TL01_CLR1_n_574, TL01_CLR1_n_575, TL01_CLR1_n_576, TL01_CLR1_n_577, TL01_CLR1_n_578 : std_logic;
  signal TL01_CLR1_n_579, TL01_CLR1_n_580, TL01_CLR1_n_581, TL01_CLR1_n_582, TL01_CLR1_n_583 : std_logic;
  signal TL01_CLR1_n_584, TL01_CLR1_n_585, TL01_CLR1_n_586, TL01_CLR1_n_587, TL01_CLR1_n_588 : std_logic;
  signal TL01_CLR1_n_589, TL01_CLR1_n_590, TL01_CLR1_n_591, TL01_CLR1_n_592, TL01_CLR1_n_593 : std_logic;
  signal TL01_CLR1_n_594, TL01_CLR1_n_595, TL01_CLR1_n_596, TL01_CLR1_n_597, TL01_CLR1_n_598 : std_logic;
  signal TL01_CLR1_n_599, TL01_CLR1_n_600, TL01_CLR1_n_601, TL01_CLR1_n_602, TL01_CLR1_n_603 : std_logic;
  signal TL01_CLR1_n_604, TL01_CLR1_n_606, TL01_CLR1_n_607, TL01_CLR1_n_608, TL01_CLR1_n_609 : std_logic;
  signal TL01_CLR1_n_610, TL01_CLR1_n_611, TL01_CLR1_n_612, TL01_CLR1_n_613, TL01_CLR1_n_614 : std_logic;
  signal TL01_CLR1_n_615, TL01_CLR1_n_616, TL01_CLR1_n_617, TL01_CLR1_n_618, TL01_CLR1_n_619 : std_logic;
  signal TL01_CLR1_n_620, TL01_CLR1_n_621, TL01_CLR1_n_622, TL01_CLR1_n_623, TL01_CLR1_n_624 : std_logic;
  signal TL01_CLR1_n_625, TL01_CLR1_n_626, TL01_CLR1_n_627, TL01_CLR1_n_628, TL01_CLR1_n_629 : std_logic;
  signal TL01_CLR1_n_630, TL01_CLR1_n_631, TL01_CLR1_n_632, TL01_CLR1_n_633, TL01_CLR1_n_634 : std_logic;
  signal TL01_CLR1_n_635, TL01_CLR1_n_636, TL01_CLR1_n_637, TL01_CLR1_n_638, TL01_CLR1_n_639 : std_logic;
  signal TL01_CLR1_n_640, TL01_CLR1_n_641, TL01_CLR1_n_642, TL01_CLR1_n_643, TL01_CLR1_n_644 : std_logic;
  signal TL01_CLR1_n_645, TL01_CLR1_n_646, TL01_CLR1_n_647, TL01_CLR1_n_648, TL01_CLR1_n_649 : std_logic;
  signal TL01_CLR1_n_650, TL01_CLR1_n_651, TL01_CLR1_n_652, TL01_CLR1_n_653, TL01_CLR1_n_654 : std_logic;
  signal TL01_CLR1_n_655, TL01_CLR1_n_656, TL01_CLR1_n_657, TL01_CLR1_n_658, TL01_CLR1_n_659 : std_logic;
  signal TL01_CLR1_n_660, TL01_CLR1_n_661, TL01_CLR1_n_662, TL01_CLR1_n_663, TL01_CLR1_n_664 : std_logic;
  signal TL01_CLR1_n_665, TL01_CLR1_n_666, TL01_CLR1_n_667, TL01_CLR1_n_668, TL01_CLR1_n_669 : std_logic;
  signal TL01_CLR1_n_670, TL01_CLR1_n_671, TL01_CLR1_n_672, TL01_CLR1_n_673, TL01_CLR1_n_674 : std_logic;
  signal TL01_CLR1_n_675, TL01_CLR1_n_676, TL01_CLR1_n_677, TL01_CLR1_n_678, TL01_CLR1_n_679 : std_logic;
  signal TL01_CLR1_n_680, TL01_CLR1_n_681, TL01_CLR1_n_682, TL01_CLR1_n_683, TL01_CLR1_n_684 : std_logic;
  signal TL01_CLR1_n_685, TL01_CLR1_n_686, TL01_CLR1_n_687, TL01_CLR1_n_688, TL01_CLR1_n_689 : std_logic;
  signal TL01_CLR1_n_690, TL01_CLR1_n_691, TL01_CLR1_n_692, TL01_CLR1_n_693, TL01_CLR1_n_694 : std_logic;
  signal TL01_CLR1_n_695, TL01_CLR1_n_696, TL01_CLR1_n_697, TL01_CLR1_n_698, TL01_CLR1_n_699 : std_logic;
  signal TL01_CLR1_n_700, TL01_CLR1_n_701, TL01_CLR1_n_702, TL01_CLR1_n_703, TL01_CLR1_n_704 : std_logic;
  signal TL01_CLR1_n_705, TL01_CLR1_n_706, TL01_CLR1_n_707, TL01_CLR1_n_708, TL01_CLR1_n_709 : std_logic;
  signal TL01_CLR1_n_710, TL01_CLR1_n_711, TL01_CLR1_n_712, TL01_CLR1_n_713, TL01_CLR1_n_714 : std_logic;
  signal TL01_CLR1_n_715, TL01_CLR1_n_716, TL01_CLR1_n_717, TL01_CLR1_n_718, TL01_CLR1_n_719 : std_logic;
  signal TL01_CLR1_n_720, TL01_CLR1_n_721, TL01_CLR1_n_722, TL01_CLR1_n_723, TL01_CLR1_n_724 : std_logic;
  signal TL01_CLR1_n_725, TL01_CLR1_n_726, TL01_CLR1_n_727, TL01_CLR1_n_728, TL01_CLR1_n_729 : std_logic;
  signal TL01_CLR1_n_730, TL01_CLR1_n_731, TL01_CLR1_n_732, TL01_CLR1_n_733, TL01_CLR1_n_734 : std_logic;
  signal TL01_CLR1_n_735, TL01_CLR1_n_736, TL01_CLR1_n_737, TL01_CLR1_n_738, TL01_CLR1_n_739 : std_logic;
  signal TL01_CLR1_n_740, TL01_CLR1_n_741, TL01_CLR1_n_742, TL01_CLR1_n_743, TL01_CLR1_n_744 : std_logic;
  signal TL01_CLR1_n_745, TL01_CLR1_n_746, TL01_CLR1_n_747, TL01_CLR1_n_748, TL01_CLR1_n_749 : std_logic;
  signal TL01_CLR1_n_750, TL01_CLR1_n_751, TL01_CLR1_n_752, TL01_CLR1_n_753, TL01_CLR1_n_754 : std_logic;
  signal TL01_CLR1_n_755, TL01_CLR1_n_756, TL01_CLR1_n_757, TL01_CLR1_n_758, TL01_CLR1_n_759 : std_logic;
  signal TL01_CLR1_n_760, TL01_CLR1_n_761, TL01_CLR1_n_762, TL01_CLR1_n_763, TL01_CLR1_n_764 : std_logic;
  signal TL01_CLR1_n_765, TL01_CLR1_n_766, TL01_CLR1_n_767, TL01_CLR1_n_768, TL01_CLR1_n_769 : std_logic;
  signal TL01_CLR1_n_770, TL01_CLR1_n_771, TL01_CLR1_n_772, TL01_CLR1_n_773, TL01_CLR1_n_774 : std_logic;
  signal TL01_CLR1_n_775, TL01_CLR1_n_776, TL01_CLR1_n_777, TL01_CLR1_n_778, TL01_CLR1_n_779 : std_logic;
  signal TL01_CLR1_n_780, TL01_CLR1_n_781, TL01_CLR1_n_782, TL01_CLR1_n_783, TL01_CLR1_n_784 : std_logic;
  signal TL01_CLR1_n_785, TL01_CLR1_n_786, TL01_CLR1_n_787, TL01_CLR1_n_788, TL01_CLR1_n_789 : std_logic;
  signal TL01_CLR1_n_790, TL01_CLR1_n_791, TL01_CLR1_n_792, TL01_CLR1_n_793, TL01_CLR1_n_794 : std_logic;
  signal TL01_CLR1_n_795, TL01_CLR1_n_796, TL01_CLR1_n_797, TL01_CLR1_n_798, TL01_CLR1_n_799 : std_logic;
  signal TL01_CLR1_n_800, TL01_CLR1_n_801, TL01_CLR1_n_802, TL01_CLR1_n_803, TL01_CLR1_n_804 : std_logic;
  signal TL01_CLR1_n_805, TL01_CLR1_n_806, TL01_CLR1_n_807, TL01_CLR1_n_808, TL01_CLR1_n_809 : std_logic;
  signal TL01_CLR1_n_810, TL01_CLR1_n_811, TL01_CLR1_n_812, TL01_CLR1_n_813, TL01_CLR1_n_814 : std_logic;
  signal TL01_CLR1_n_815, TL01_CLR1_n_816, TL01_CLR1_n_817, TL01_CLR1_n_818, TL01_CLR1_n_819 : std_logic;
  signal TL01_CLR1_n_820, TL01_CLR1_n_821, TL01_CLR1_n_822, TL01_CLR1_n_823, TL01_CLR1_n_824 : std_logic;
  signal TL01_CLR1_n_825, TL01_CLR1_n_826, TL01_CLR1_n_827, TL01_CLR1_n_828, TL01_CLR1_n_829 : std_logic;
  signal TL01_CLR1_n_830, TL01_CLR1_n_831, TL01_CLR1_n_832, TL01_CLR1_n_833, TL01_CLR1_n_834 : std_logic;
  signal TL01_CLR1_n_835, TL01_CLR1_n_836, TL01_CLR1_n_837, TL01_CLR1_n_838, TL01_CLR1_n_839 : std_logic;
  signal TL01_CLR1_n_840, TL01_CLR1_n_841, TL01_CLR1_n_842, TL01_CLR1_n_843, TL01_CLR1_n_844 : std_logic;
  signal TL01_CLR1_n_845, TL01_CLR1_n_846, TL01_CLR1_n_847, TL01_CLR1_n_848, TL01_CLR1_n_849 : std_logic;
  signal TL01_CLR1_n_850, TL01_CLR1_n_851, TL01_CLR1_n_852, TL01_CLR1_n_853, TL01_CLR1_n_854 : std_logic;
  signal TL01_CLR1_n_855, TL01_CLR1_n_856, TL01_CLR1_n_857, TL01_CLR1_n_858, TL01_CLR1_n_859 : std_logic;
  signal TL01_CLR1_n_860, TL01_CLR1_n_861, TL01_CLR1_n_862, TL01_CLR1_n_863, TL01_CLR1_n_864 : std_logic;
  signal TL01_CLR1_n_865, TL01_CLR1_n_866, TL01_CLR1_n_867, TL01_CLR1_n_868, TL01_CLR1_n_869 : std_logic;
  signal TL01_CLR1_n_870, TL01_CLR1_n_871, TL01_CLR1_n_872, TL01_CLR1_n_873, TL01_CLR1_n_874 : std_logic;
  signal TL01_CLR1_n_875, TL01_CLR1_n_876, TL01_CLR1_n_877, TL01_CLR1_n_878, TL01_CLR1_n_879 : std_logic;
  signal TL01_CLR1_n_880, TL01_CLR1_n_881, TL01_CLR1_n_882, TL01_CLR1_n_883, TL01_CLR1_n_884 : std_logic;
  signal TL01_CLR1_n_885, TL01_CLR1_n_886, TL01_CLR1_n_887, TL01_CLR1_n_888, TL01_CLR1_n_889 : std_logic;
  signal TL01_CLR1_n_890, TL01_CLR1_n_891, TL01_CLR1_n_892, TL01_CLR1_n_893, TL01_CLR1_n_894 : std_logic;
  signal TL01_CLR1_n_895, TL01_CLR1_n_896, TL01_CLR1_n_897, TL01_CLR1_n_898, TL01_CLR1_n_899 : std_logic;
  signal TL01_CLR1_n_900, TL01_CLR1_n_901, TL01_CLR1_n_902, TL01_CLR1_n_903, TL01_CLR1_n_904 : std_logic;
  signal TL01_CLR1_n_905, TL01_CLR1_n_906, TL01_CLR1_n_907, TL01_CLR1_n_908, TL01_CLR1_n_909 : std_logic;
  signal TL01_CLR1_n_910, TL01_CLR1_n_911, TL01_CLR1_n_912, TL01_CLR1_n_913, TL01_CLR1_n_914 : std_logic;
  signal TL01_CLR1_n_915, TL01_CLR1_n_916, TL01_CLR1_n_917, TL01_CLR1_n_918, TL01_CLR1_n_919 : std_logic;
  signal TL01_CLR1_n_920, TL01_CLR1_n_921, TL01_CLR1_n_922, TL01_CLR1_n_923, TL01_CLR1_n_924 : std_logic;
  signal TL01_CLR1_n_925, TL01_CLR1_n_926, TL01_CLR1_n_927, TL01_CLR1_n_928, TL01_CLR1_n_929 : std_logic;
  signal TL01_CLR1_n_930, TL01_CLR1_n_931, TL01_CLR1_n_932, TL01_CLR1_n_933, TL01_CLR1_n_934 : std_logic;
  signal TL01_CLR1_n_935, TL01_CLR1_n_936, TL01_CLR1_n_937, TL01_CLR1_n_938, TL01_CLR1_n_939 : std_logic;
  signal TL01_CLR1_n_940, TL01_CLR1_n_941, TL01_CLR1_n_942, TL01_CLR1_n_943, TL01_CLR1_n_944 : std_logic;
  signal TL01_CLR1_n_945, TL01_CLR1_n_946, TL01_CLR1_n_947, TL01_CLR1_n_948, TL01_CLR1_n_949 : std_logic;
  signal TL01_CLR1_n_950, TL01_CLR1_n_951, TL01_CLR1_n_952, TL01_CLR1_n_953, TL01_CLR1_n_954 : std_logic;
  signal TL01_CLR1_n_955, TL01_CLR1_n_956, TL01_CLR1_n_957, TL01_CLR1_n_958, TL01_CLR1_n_959 : std_logic;
  signal TL01_CLR1_n_960, TL01_CLR1_n_961, TL01_CLR1_n_962, TL01_CLR1_n_963, TL01_CLR1_n_964 : std_logic;
  signal TL01_CLR1_n_965, TL01_CLR1_n_966, TL01_CLR1_n_967, TL01_CLR1_n_968, TL01_CLR1_n_969 : std_logic;
  signal TL01_CLR1_n_970, TL01_CLR1_n_971, TL01_CLR1_n_972, TL01_CLR1_n_973, TL01_CLR1_n_974 : std_logic;
  signal TL01_CLR1_n_975, TL01_CLR1_n_976, TL01_CLR1_n_977, TL01_CLR1_n_978, TL01_CLR1_n_979 : std_logic;
  signal TL01_CLR1_n_980, TL01_CLR1_n_981, TL01_CLR1_n_982, TL01_CLR1_n_983, TL01_CLR1_n_984 : std_logic;
  signal TL01_CLR1_n_985, TL01_CLR1_n_986, TL01_CLR1_n_987, TL01_CLR1_n_988, TL01_CLR1_n_989 : std_logic;
  signal TL01_CLR1_n_990, TL01_CLR1_n_991, TL01_CLR1_n_992, TL01_CLR1_n_993, TL01_CLR1_n_994 : std_logic;
  signal TL01_CLR1_n_995, TL01_CLR1_n_996, TL01_CLR1_n_997, TL01_CLR1_n_998, TL01_CLR1_n_999 : std_logic;
  signal TL01_CLR1_n_1000, TL01_CLR1_n_1001, TL01_CLR1_n_1002, TL01_CLR1_n_1003, TL01_CLR1_n_1004 : std_logic;
  signal TL01_CLR1_n_1005, TL01_CLR1_n_1006, TL01_CLR1_n_1007, TL01_CLR1_n_1008, TL01_CLR1_n_1009 : std_logic;
  signal TL01_CLR1_n_1010, TL01_CLR1_n_1011, TL01_CLR1_n_1012, TL01_CLR1_n_1013, TL01_CLR1_n_1014 : std_logic;
  signal TL01_CLR1_n_1015, TL01_CLR1_n_1016, TL01_CLR1_n_1017, TL01_CLR1_n_1018, TL01_CLR1_n_1019 : std_logic;
  signal TL01_CLR1_n_1020, TL01_CLR1_n_1021, TL01_CLR1_n_1022, TL01_CLR1_n_1023, TL01_CLR1_n_1024 : std_logic;
  signal TL01_CLR1_n_1025, TL01_CLR1_n_1026, TL01_CLR1_n_1027, TL01_CLR1_n_1028, TL01_CLR1_n_1029 : std_logic;
  signal TL01_CLR1_n_1030, TL01_CLR1_n_1031, TL01_CLR1_n_1032, TL01_CLR1_n_1033, TL01_CLR1_n_1034 : std_logic;
  signal TL01_CLR1_n_1035, TL01_CLR1_n_1036, TL01_CLR1_n_1037, TL01_CLR1_n_1038, TL01_CLR1_n_1039 : std_logic;
  signal TL01_CLR1_n_1040, TL01_CLR1_n_1041, TL01_CLR1_n_1042, TL01_CLR1_n_1043, TL01_CLR1_n_1044 : std_logic;
  signal TL01_CLR1_n_1045, TL01_CLR1_n_1046, TL01_CLR1_n_1047, TL01_CLR1_n_1048, TL01_CLR1_n_1049 : std_logic;
  signal TL01_CLR1_n_1050, TL01_CLR1_n_1051, TL01_CLR1_n_1052, TL01_CLR1_n_1053, TL01_CLR1_n_1054 : std_logic;
  signal TL01_CLR1_n_1055, TL01_CLR1_n_1056, TL01_CLR1_n_1057, TL01_CLR1_n_1058, TL01_CLR1_n_1059 : std_logic;
  signal TL01_CLR1_n_1060, TL01_CLR1_n_1061, TL01_CLR1_n_1062, TL01_CLR1_n_1063, TL01_CLR1_n_1064 : std_logic;
  signal TL01_CLR1_n_1065, TL01_CLR1_n_1066, TL01_CLR1_n_1067, TL01_CLR1_n_1068, TL01_CLR1_n_1069 : std_logic;
  signal TL01_CLR1_n_1070, TL01_CLR1_n_1071, TL01_CLR1_n_1072, TL01_CLR1_n_1073, TL01_CLR1_n_1074 : std_logic;
  signal TL01_CLR1_n_1075, TL01_CLR1_n_1076, TL01_CLR1_n_1077, TL01_CLR1_n_1078, TL01_CLR1_n_1079 : std_logic;
  signal TL01_CLR1_n_1080, TL01_CLR1_n_1081, TL01_CLR1_n_1082, TL01_CLR1_n_1083, TL01_CLR1_n_1084 : std_logic;
  signal TL01_CLR1_n_1085, TL01_CLR1_n_1086, TL01_CLR1_n_1087, TL01_CLR1_n_1088, TL01_CLR1_n_1089 : std_logic;
  signal TL01_CLR1_n_1090, TL01_CLR1_n_1091, TL01_CLR1_n_1092, TL01_CLR1_n_1093, TL01_CLR1_n_1094 : std_logic;
  signal TL01_CLR1_n_1095, TL01_CLR1_n_1096, TL01_CLR1_n_1097, TL01_CLR1_n_1098, TL01_CLR1_n_1099 : std_logic;
  signal TL01_CLR1_n_1100, TL01_CLR1_n_1101, TL01_CLR1_n_1102, TL01_CLR1_n_1103, TL01_CLR1_n_1104 : std_logic;
  signal TL01_CLR1_n_1105, TL01_CLR1_n_1106, TL01_CLR1_n_1107, TL01_CLR1_n_1108, TL01_CLR1_n_1109 : std_logic;
  signal TL01_CLR1_n_1110, TL01_CLR1_n_1111, TL01_CLR1_n_1112, TL01_CLR1_n_1113, TL01_CLR1_n_1114 : std_logic;
  signal TL01_CLR1_n_1115, TL01_CLR1_n_1116, TL01_CLR1_n_1117, TL01_CLR1_n_1118, TL01_CLR1_n_1119 : std_logic;
  signal TL01_CLR1_n_1120, TL01_CLR1_n_1121, TL01_CLR1_n_1122, TL01_CLR1_n_1123, TL01_CLR1_n_1124 : std_logic;
  signal TL01_CLR1_n_1125, TL01_CLR1_n_1126, TL01_CLR1_n_1127, TL01_CLR1_n_1128, TL01_CLR1_n_1129 : std_logic;
  signal TL01_CLR1_n_1130, TL01_CLR1_n_1131, TL01_CLR1_n_1132, TL01_CLR1_n_1133, TL01_CLR1_n_1134 : std_logic;
  signal TL01_CLR1_n_1135, TL01_CLR1_n_1136, TL01_CLR1_n_1137, TL01_CLR1_n_1138, TL01_CLR1_n_1139 : std_logic;
  signal TL01_CLR1_n_1140, TL01_CLR1_n_1141, TL01_CLR1_n_1142, TL01_CLR1_n_1143, TL01_CLR1_n_1144 : std_logic;
  signal TL01_CLR1_n_1145, TL01_CLR1_n_1146, TL01_CLR1_n_1147, TL01_CLR1_n_1148, TL01_CLR1_n_1149 : std_logic;
  signal TL01_CLR1_n_1150, TL01_CLR1_n_1151, TL01_CLR1_n_1152, TL01_CLR1_n_1153, TL01_CLR1_n_1154 : std_logic;
  signal TL01_CLR1_n_1155, TL01_CLR1_n_1156, TL01_CLR1_n_1157, TL01_CLR1_n_1158, TL01_CLR1_n_1159 : std_logic;
  signal TL01_CLR1_n_1160, TL01_CLR1_n_1161, TL01_CLR1_n_1162, TL01_CLR1_n_1163, TL01_CLR1_n_1164 : std_logic;
  signal TL01_CLR1_n_1165, TL01_CLR1_n_1166, TL01_CLR1_n_1167, TL01_CLR1_n_1168, TL01_CLR1_n_1169 : std_logic;
  signal TL01_CLR1_n_1170, TL01_CLR1_n_1171, TL01_CLR1_n_1172, TL01_CLR1_n_1173, TL01_CLR1_n_1174 : std_logic;
  signal TL01_CLR1_n_1175, TL01_CLR1_n_1176, TL01_CLR1_n_1177, TL01_CLR1_n_1178, TL01_CLR1_n_1179 : std_logic;
  signal TL01_CLR1_n_1180, TL01_CLR1_n_1181, TL01_CLR1_n_1182, TL01_CLR1_n_1183, TL01_CLR1_n_1184 : std_logic;
  signal TL01_CLR1_n_1185, TL01_CLR1_n_1186, TL01_CLR1_n_1187, TL01_CLR1_n_1188, TL01_CLR1_n_1189 : std_logic;
  signal TL01_CLR1_n_1190, TL01_CLR1_n_1191, TL01_CLR1_n_1192, TL01_CLR1_n_1193, TL01_CLR1_n_1194 : std_logic;
  signal TL01_CLR1_n_1195, TL01_CLR1_n_1196, TL01_CLR1_n_1197, TL01_CLR1_n_1198, TL01_CLR1_n_1199 : std_logic;
  signal TL01_CLR1_n_1200, TL01_CLR1_n_1201, TL01_CLR1_n_1202, TL01_CLR1_n_1203, TL01_CLR1_n_1204 : std_logic;
  signal TL01_CLR1_n_1205, TL01_CLR1_n_1206, TL01_CLR1_n_1207, TL01_CLR1_n_1208, TL01_CLR1_n_1209 : std_logic;
  signal TL01_CLR1_n_1210, TL01_CLR1_n_1211, TL01_CLR1_n_1212, TL01_CLR1_n_1213, TL01_CLR1_n_1214 : std_logic;
  signal TL01_CLR1_n_1215, TL01_CLR1_n_1216, TL01_CLR1_n_1217, TL01_CLR1_n_1218, TL01_CLR1_n_1219 : std_logic;
  signal TL01_CLR1_n_1220, TL01_CLR1_n_1221, TL01_CLR1_n_1222, TL01_CLR1_n_1223, TL01_CLR1_n_1224 : std_logic;
  signal TL01_CLR1_n_1225, TL01_CLR1_n_1226, TL01_CLR1_n_1227, TL01_CLR1_n_1228, TL01_CLR1_n_1229 : std_logic;
  signal TL01_CLR1_n_1230, TL01_CLR1_n_1231, TL01_CLR1_n_1232, TL01_CLR1_n_1233, TL01_CLR1_n_1234 : std_logic;
  signal TL01_CLR1_n_1235, TL01_CLR1_n_1236, TL01_CLR1_n_1237, TL01_CLR1_n_1238, TL01_CLR1_n_1239 : std_logic;
  signal TL01_CLR1_n_1240, TL01_CLR1_n_1241, TL01_CLR1_n_1242, TL01_CLR1_n_1243, TL01_CLR1_n_1244 : std_logic;
  signal TL01_CLR1_n_1245, TL01_CLR1_n_1246, TL01_CLR1_n_1247, TL01_CLR1_n_1248, TL01_CLR1_n_1249 : std_logic;
  signal TL01_CLR1_n_1250, TL01_CLR1_n_1251, TL01_CLR1_n_1252, TL01_CLR1_n_1253, TL01_CLR1_n_1254 : std_logic;
  signal TL01_CLR1_n_1255, TL01_CLR1_n_1256, TL01_CLR1_n_1257, TL01_CLR1_n_1258, TL01_CLR1_n_1259 : std_logic;
  signal TL01_CLR1_n_1260, TL01_CLR1_n_1261, TL01_CLR1_n_1262, TL01_CLR1_n_1263, TL01_CLR1_n_1264 : std_logic;
  signal TL01_CLR1_n_1265, TL01_CLR1_n_1266, TL01_CLR1_n_1267, TL01_CLR1_n_1268, TL01_CLR1_n_1269 : std_logic;
  signal TL01_CLR1_n_1270, TL01_CLR1_n_1271, TL01_CLR1_n_1272, TL01_CLR1_n_1273, TL01_CLR1_n_1274 : std_logic;
  signal TL01_CLR1_n_1275, TL01_CLR1_n_1276, TL01_CLR1_n_1277, TL01_CLR1_n_1278, TL01_CLR1_n_1279 : std_logic;
  signal TL01_CLR1_n_1280, TL01_CLR1_n_1281, TL01_CLR1_n_1282, TL01_CLR1_n_1283, TL01_CLR1_n_1284 : std_logic;
  signal TL01_CLR1_n_1285, TL01_CLR1_n_1286, TL01_CLR1_n_1287, TL01_CLR1_n_1288, TL01_CLR1_n_1289 : std_logic;
  signal TL01_CLR1_n_1290, TL01_CLR1_n_1291, TL01_CLR1_n_1292, TL01_CLR1_n_1293, TL01_CLR1_n_1294 : std_logic;
  signal TL01_CLR1_n_1295, TL01_CLR1_n_1296, TL01_CLR1_n_1297, TL01_CLR1_n_1298, TL01_CLR1_n_1299 : std_logic;
  signal TL01_CLR1_n_1300, TL01_CLR1_n_1301, TL01_CLR1_n_1302, TL01_CLR1_n_1303, TL01_CLR1_n_1304 : std_logic;
  signal TL01_CLR1_n_1305, TL01_CLR1_n_1306, TL01_CLR1_n_1307, TL01_CLR1_n_1308, TL01_CLR1_n_1309 : std_logic;
  signal TL01_CLR1_n_1310, TL01_CLR1_n_1311, TL01_CLR1_n_1312, TL01_CLR1_n_1313, TL01_CLR1_n_1314 : std_logic;
  signal TL01_CLR1_n_1315, TL01_CLR1_n_1316, TL01_CLR1_n_1317, TL01_CLR1_n_1318, TL01_CLR1_n_1319 : std_logic;
  signal TL01_CLR1_n_1320, TL01_CLR1_n_1321, TL01_CLR1_n_1322, TL01_CLR1_n_1323, TL01_CLR1_n_1324 : std_logic;
  signal TL01_CLR1_n_1325, TL01_CLR1_n_1326, TL01_CLR1_n_1327, TL01_CLR1_n_1328, TL01_CLR1_n_1329 : std_logic;
  signal TL01_CLR1_n_1330, TL01_CLR1_n_1331, TL01_CLR1_n_1332, TL01_CLR1_n_1333, TL01_CLR1_n_1334 : std_logic;
  signal TL01_CLR1_n_1335, TL01_CLR1_n_1336, TL01_CLR1_n_1337, TL01_CLR1_n_1338, TL01_CLR1_n_1339 : std_logic;
  signal TL01_CLR1_n_1340, TL01_CLR1_n_1341, TL01_CLR1_n_1342, TL01_CLR1_n_1343, TL01_CLR1_n_1344 : std_logic;
  signal TL01_CLR1_n_1345, TL01_CLR1_n_1346, TL01_CLR1_n_1347, TL01_CLR1_n_1348, TL01_CLR1_n_1349 : std_logic;
  signal TL01_CLR1_n_1350, TL01_CLR1_n_1351, TL01_CLR1_n_1352, TL01_CLR1_n_1353, TL01_CLR1_n_1354 : std_logic;
  signal TL01_CLR1_n_1355, TL01_CLR1_n_1356, TL01_CLR1_n_1357, TL01_CLR1_n_1358, TL01_CLR1_n_1359 : std_logic;
  signal TL01_CLR1_n_1360, TL01_CLR1_n_1361, TL01_CLR1_n_1362, TL01_CLR1_n_1363, TL01_CLR1_n_1364 : std_logic;
  signal TL01_CLR1_n_1365, TL01_CLR1_n_1366, TL01_CLR1_n_1367, TL01_CLR1_n_1368, TL01_CLR1_n_1369 : std_logic;
  signal TL01_CLR1_n_1370, TL01_CLR1_n_1371, TL01_CLR1_n_1372, TL01_CLR1_n_1373, TL01_CLR1_n_1374 : std_logic;
  signal TL01_CLR1_n_1375, TL01_CLR1_n_1376, TL01_CLR1_n_1377, TL01_CLR1_n_1378, TL01_CLR1_n_1379 : std_logic;
  signal TL01_CLR1_n_1380, TL01_CLR1_n_1381, TL01_CLR1_n_1382, TL01_CLR1_n_1383, TL01_CLR1_n_1384 : std_logic;
  signal TL01_CLR1_n_1385, TL01_CLR1_n_1386, TL01_CLR1_n_1387, TL01_CLR1_n_1388, TL01_CLR1_n_1389 : std_logic;
  signal TL01_CLR1_n_1390, TL01_CLR1_n_1391, TL01_CLR1_n_1392, TL01_CLR1_n_1393, TL01_CLR1_n_1394 : std_logic;
  signal TL01_CLR1_n_1395, TL01_CLR1_n_1396, TL01_CLR1_n_1397, TL01_CLR1_n_1398, TL01_CLR1_n_1399 : std_logic;
  signal TL01_CLR1_n_1400, TL01_CLR1_n_1401, TL01_CLR1_n_1402, TL01_CLR1_n_1403, TL01_CLR1_n_1404 : std_logic;
  signal TL01_CLR1_n_1405, TL01_CLR1_n_1406, TL01_CLR1_n_1407, TL01_CLR1_n_1408, TL01_CLR1_n_1409 : std_logic;
  signal TL01_CLR1_n_1410, TL01_CLR1_n_1411, TL01_CLR1_n_1412, TL01_CLR1_n_1413, TL01_CLR1_n_1414 : std_logic;
  signal TL01_CLR1_n_1415, TL01_CLR1_n_1416, TL01_CLR1_n_1417, TL01_CLR1_n_1418, TL01_CLR1_n_1419 : std_logic;
  signal TL01_CLR1_n_1420, TL01_CLR1_n_1421, TL01_CLR1_n_1422, TL01_CLR1_n_1423, TL01_CLR1_n_1424 : std_logic;
  signal TL01_CLR1_n_1425, TL01_CLR1_n_1426, TL01_CLR1_n_1427, TL01_CLR1_n_1428, TL01_CLR1_n_1429 : std_logic;
  signal TL01_CLR1_n_1430, TL01_CLR1_n_1431, TL01_CLR1_n_1432, TL01_CLR1_n_1433, TL01_CLR1_n_1434 : std_logic;
  signal TL01_CLR1_n_1435, TL01_CLR1_n_1436, TL01_CLR1_n_1437, TL01_CLR1_n_1438, TL01_CLR1_n_1439 : std_logic;
  signal TL01_CLR1_n_1440, TL01_CLR1_n_1441, TL01_CLR1_n_1442, TL01_CLR1_n_1443, TL01_CLR1_n_1444 : std_logic;
  signal TL01_CLR1_n_1445, TL01_CLR1_n_1446, TL01_CLR1_n_1447, TL01_CLR1_n_1448, TL01_CLR1_n_1449 : std_logic;
  signal TL01_CLR1_n_1450, TL01_CLR1_n_1451, TL01_CLR1_n_1452, TL01_CLR1_n_1453, TL01_CLR1_n_1454 : std_logic;
  signal TL01_CLR1_n_1455, TL01_CLR1_n_1456, TL01_CLR1_n_1457, TL01_CLR1_n_1458, TL01_CLR1_n_1459 : std_logic;
  signal TL01_CLR1_n_1460, TL01_CLR1_n_1461, TL01_CLR1_n_1462, TL01_CLR1_n_1463, TL01_CLR1_n_1464 : std_logic;
  signal TL01_CLR1_n_1465, TL01_CLR1_n_1466, TL01_CLR1_n_1467, TL01_CLR1_n_1468, TL01_CLR1_n_1469 : std_logic;
  signal TL01_CLR1_n_1470, TL01_CLR1_n_1471, TL01_CLR1_n_1472, TL01_CLR1_n_1473, TL01_CLR1_n_1475 : std_logic;
  signal TL01_CLR1_n_1477, TL01_CLR1_n_1478, TL01_CLR1_n_1479, TL01_CLR1_n_1480, TL01_CLR1_n_1481 : std_logic;
  signal TL01_CLR1_n_1482, TL01_CLR1_n_1483, TL01_CLR1_n_1484, TL01_CLR1_n_1486, TL01_CLR1_n_1487 : std_logic;
  signal TL01_CLR1_n_1488, TL01_CLR1_n_1489, TL01_CLR1_n_1490, TL01_CLR1_n_1491, TL01_CLR1_n_1492 : std_logic;
  signal TL01_CLR1_n_1493, TL01_CLR1_n_1494, TL01_CLR1_n_1495, TL01_CLR1_n_1561, TL01_CLR1_n_1562 : std_logic;
  signal TL01_CLR1_n_1563, TL01_CLR1_n_1564, TL01_CLR1_n_1565, TL01_SCNR1_hcount_reset, TL01_SCNR1_vcount_reset : std_logic;
  signal TL01_n_0, TL01_n_1, TL01_n_2, TL01_n_3, TL01_n_4 : std_logic;
  signal TL01_n_5, TL01_n_6, TL01_n_7, TL01_n_8, TL01_n_9 : std_logic;
  signal TL01_n_10, TL01_n_11, TL01_n_12, TL01_n_13, TL01_n_14 : std_logic;
  signal TL01_n_15, TL01_n_16, TL01_n_17, TL01_n_18, TL01_n_19 : std_logic;
  signal TL01_n_20, TL01_n_21, TL01_n_22, TL01_n_23, TL01_n_24 : std_logic;
  signal TL01_n_25, TL01_n_26, TL01_n_27, TL01_n_28, TL01_n_29 : std_logic;
  signal TL01_n_30, TL01_n_31, TL01_n_32, TL01_n_33, TL01_n_34 : std_logic;
  signal TL01_n_35, TL01_n_36, TL01_n_37, TL01_n_38, TL01_n_39 : std_logic;
  signal TL01_n_40, TL01_n_41, TL01_n_42, TL01_n_43, TL01_n_44 : std_logic;
  signal TL01_n_45, TL01_n_46, TL01_n_47, TL01_n_48, TL01_n_49 : std_logic;
  signal TL01_n_50, TL01_n_51, TL01_n_52, TL01_n_53, TL01_n_54 : std_logic;
  signal TL01_n_55, TL01_n_56, TL01_n_57, TL01_n_58, TL01_n_59 : std_logic;
  signal TL01_n_60, TL01_n_61, TL01_n_62, TL01_n_63, TL02_PHS0_sel_0 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_1, TL02_PHS1_knockback_mul_35_64_n_2, TL02_PHS1_knockback_mul_35_64_n_3, TL02_PHS1_knockback_mul_35_64_n_4, TL02_PHS1_knockback_mul_35_64_n_5 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_6, TL02_PHS1_knockback_mul_35_64_n_7, TL02_PHS1_knockback_mul_35_64_n_8, TL02_PHS1_knockback_mul_35_64_n_9, TL02_PHS1_knockback_mul_35_64_n_10 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_11, TL02_PHS1_knockback_mul_35_64_n_12, TL02_PHS1_knockback_mul_35_64_n_13, TL02_PHS1_knockback_mul_35_64_n_14, TL02_PHS1_knockback_mul_35_64_n_15 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_16, TL02_PHS1_knockback_mul_35_64_n_17, TL02_PHS1_knockback_mul_35_64_n_18, TL02_PHS1_knockback_mul_35_64_n_19, TL02_PHS1_knockback_mul_35_64_n_20 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_21, TL02_PHS1_knockback_mul_35_64_n_22, TL02_PHS1_knockback_mul_35_64_n_23, TL02_PHS1_knockback_mul_35_64_n_24, TL02_PHS1_knockback_mul_35_64_n_25 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_26, TL02_PHS1_knockback_mul_35_64_n_27, TL02_PHS1_knockback_mul_35_64_n_28, TL02_PHS1_knockback_mul_35_64_n_29, TL02_PHS1_knockback_mul_35_64_n_30 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_31, TL02_PHS1_knockback_mul_35_64_n_32, TL02_PHS1_knockback_mul_35_64_n_33, TL02_PHS1_knockback_mul_35_64_n_34, TL02_PHS1_knockback_mul_35_64_n_35 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_36, TL02_PHS1_knockback_mul_35_64_n_37, TL02_PHS1_knockback_mul_35_64_n_38, TL02_PHS1_knockback_mul_35_64_n_39, TL02_PHS1_knockback_mul_35_64_n_40 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_41, TL02_PHS1_knockback_mul_35_64_n_42, TL02_PHS1_knockback_mul_35_64_n_43, TL02_PHS1_knockback_mul_35_64_n_44, TL02_PHS1_knockback_mul_35_64_n_45 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_46, TL02_PHS1_knockback_mul_35_64_n_47, TL02_PHS1_knockback_mul_35_64_n_48, TL02_PHS1_knockback_mul_35_64_n_49, TL02_PHS1_knockback_mul_35_64_n_50 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_51, TL02_PHS1_knockback_mul_35_64_n_52, TL02_PHS1_knockback_mul_35_64_n_53, TL02_PHS1_knockback_mul_35_64_n_54, TL02_PHS1_knockback_mul_35_64_n_55 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_56, TL02_PHS1_knockback_mul_35_64_n_57, TL02_PHS1_knockback_mul_35_64_n_58, TL02_PHS1_knockback_mul_35_64_n_59, TL02_PHS1_knockback_mul_35_64_n_60 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_62, TL02_PHS1_knockback_mul_35_64_n_63, TL02_PHS1_knockback_mul_35_64_n_64, TL02_PHS1_knockback_mul_35_64_n_65, TL02_PHS1_knockback_mul_35_64_n_66 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_67, TL02_PHS1_knockback_mul_35_64_n_68, TL02_PHS1_knockback_mul_35_64_n_69, TL02_PHS1_knockback_mul_35_64_n_70, TL02_PHS1_knockback_mul_35_64_n_71 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_72, TL02_PHS1_knockback_mul_35_64_n_73, TL02_PHS1_knockback_mul_35_64_n_74, TL02_PHS1_knockback_mul_35_64_n_75, TL02_PHS1_knockback_mul_35_64_n_76 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_77, TL02_PHS1_knockback_mul_35_64_n_78, TL02_PHS1_knockback_mul_35_64_n_79, TL02_PHS1_knockback_mul_35_64_n_80, TL02_PHS1_knockback_mul_35_64_n_81 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_82, TL02_PHS1_knockback_mul_35_64_n_83, TL02_PHS1_knockback_mul_35_64_n_84, TL02_PHS1_knockback_mul_35_64_n_85, TL02_PHS1_knockback_mul_35_64_n_86 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_87, TL02_PHS1_knockback_mul_35_64_n_89, TL02_PHS1_knockback_mul_35_64_n_90, TL02_PHS1_knockback_mul_35_64_n_91, TL02_PHS1_knockback_mul_35_64_n_92 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_93, TL02_PHS1_knockback_mul_35_64_n_94, TL02_PHS1_knockback_mul_35_64_n_95, TL02_PHS1_knockback_mul_35_64_n_96, TL02_PHS1_knockback_mul_35_64_n_97 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_98, TL02_PHS1_knockback_mul_35_64_n_99, TL02_PHS1_knockback_mul_35_64_n_100, TL02_PHS1_knockback_mul_35_64_n_101, TL02_PHS1_knockback_mul_35_64_n_102 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_103, TL02_PHS1_knockback_mul_35_64_n_104, TL02_PHS1_knockback_mul_35_64_n_105, TL02_PHS1_knockback_mul_35_64_n_106, TL02_PHS1_knockback_mul_35_64_n_107 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_108, TL02_PHS1_knockback_mul_35_64_n_109, TL02_PHS1_knockback_mul_35_64_n_110, TL02_PHS1_knockback_mul_35_64_n_111, TL02_PHS1_knockback_mul_35_64_n_112 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_113, TL02_PHS1_knockback_mul_35_64_n_114, TL02_PHS1_knockback_mul_35_64_n_115, TL02_PHS1_knockback_mul_35_64_n_116, TL02_PHS1_knockback_mul_35_64_n_117 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_119, TL02_PHS1_knockback_mul_35_64_n_120, TL02_PHS1_knockback_mul_35_64_n_121, TL02_PHS1_knockback_mul_35_64_n_122, TL02_PHS1_knockback_mul_35_64_n_123 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_124, TL02_PHS1_knockback_mul_35_64_n_125, TL02_PHS1_knockback_mul_35_64_n_126, TL02_PHS1_knockback_mul_35_64_n_127, TL02_PHS1_knockback_mul_35_64_n_128 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_129, TL02_PHS1_knockback_mul_35_64_n_130, TL02_PHS1_knockback_mul_35_64_n_131, TL02_PHS1_knockback_mul_35_64_n_132, TL02_PHS1_knockback_mul_35_64_n_134 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_135, TL02_PHS1_knockback_mul_35_64_n_136, TL02_PHS1_knockback_mul_35_64_n_137, TL02_PHS1_knockback_mul_35_64_n_138, TL02_PHS1_knockback_mul_35_64_n_139 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_141, TL02_PHS1_knockback_mul_35_64_n_142, TL02_PHS1_knockback_mul_35_64_n_143, TL02_PHS1_knockback_mul_35_64_n_144, TL02_PHS1_knockback_mul_35_64_n_145 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_146, TL02_PHS1_knockback_mul_35_64_n_147, TL02_PHS1_knockback_mul_35_64_n_148, TL02_PHS1_knockback_mul_35_64_n_149, TL02_PHS1_knockback_mul_35_64_n_150 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_151, TL02_PHS1_knockback_mul_35_64_n_152, TL02_PHS1_knockback_mul_35_64_n_153, TL02_PHS1_knockback_mul_35_64_n_154, TL02_PHS1_knockback_mul_35_64_n_155 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_156, TL02_PHS1_knockback_mul_35_64_n_157, TL02_PHS1_knockback_mul_35_64_n_158, TL02_PHS1_knockback_mul_35_64_n_160, TL02_PHS1_knockback_mul_35_64_n_162 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_164, TL02_PHS1_knockback_mul_35_64_n_166, TL02_PHS1_knockback_mul_35_64_n_168, TL02_PHS1_knockback_mul_35_64_n_171, TL02_PHS1_knockback_mul_35_64_n_173 : std_logic;
  signal TL02_PHS1_knockback_mul_35_64_n_199, TL02_PHS1_knockback_mul_35_64_n_200, TL02_PHS1_knockback_mul_35_64_n_201, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_6, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_7, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_8 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_9, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_10, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_11, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_12, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_13 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_14, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_15, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_16, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_17, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_18 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_19, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_20, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_21, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_22, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_23 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_24, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_25, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_26, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_27, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_28 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_29, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_30, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_31, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_32, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_33 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_34, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_35, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_36, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_37, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_38 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_39, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_40, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_41, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_42, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_43 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_44, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_45, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_46, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_47, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_48 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_49, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_50, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_51, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_52, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_53 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_54, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_55, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_56, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_57, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_58 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_59, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_60, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_62, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_63, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_64 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_65, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_66, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_67, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_68, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_69 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_70, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_71, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_72, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_73, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_74 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_75, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_76, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_77, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_78, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_79 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_80, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_81, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_82, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_83, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_84 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_85, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_86, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_87, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_89, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_90 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_91, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_92, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_93, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_94, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_95 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_96, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_97, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_98, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_99, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_100 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_101, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_102, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_103, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_104, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_105 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_106, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_107, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_108, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_109, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_110 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_111, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_112, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_113, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_114, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_115 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_116, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_117, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_119, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_120, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_121 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_122, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_123, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_124, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_125, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_126 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_127, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_128, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_129, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_130, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_131 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_132, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_134, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_135, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_136, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_137 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_138, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_139, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_141, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_142, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_143 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_144, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_145, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_146, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_147, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_148 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_149, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_150, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_151, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_152, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_153 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_154, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_155, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_156, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_157, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_158 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_160, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_162, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_164, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_166, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_168 : std_logic;
  signal TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_171, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_173, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_199, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_200, TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_201 : std_logic;
  signal TL02_kb_y_0, TL02_kb_y_1, TL02_kb_y_2, TL02_kb_y_3, TL02_kb_y_4 : std_logic;
  signal TL02_kb_y_5, TL02_kb_y_6, TL02_n_438, TL02_n_439, TL02_n_440 : std_logic;
  signal TL02_n_441, TL02_n_442, TL02_n_443, TL02_n_444, TL02_n_445 : std_logic;
  signal TL02_n_446, TL02_n_447, TL02_n_448, TL02_n_449, TL02_n_450 : std_logic;
  signal TL02_n_451, TL02_n_452, TL02_n_453, TL02_n_454, TL02_n_456 : std_logic;
  signal TL02_n_457, TL02_n_458, TL02_n_459, TL02_n_460, TL02_n_461 : std_logic;
  signal TL02_n_462, TL02_n_463, TL02_n_592, TL02_n_594, TL02_n_595 : std_logic;
  signal TL02_n_596, TL02_n_597, TL02_n_598, TL02_n_599, TL02_n_600 : std_logic;
  signal TL02_n_601, TL04_count_reset, TL04_des_clk_buffered, TL04_driver_pulse_count_0, TL04_driver_pulse_count_1 : std_logic;
  signal TL04_driver_pulse_count_2, TL04_driver_state_0, TL04_driver_state_1, TL04_driver_state_2, TL04_jump_button_p1 : std_logic;
  signal TL04_jump_button_p2, TL04_jump_p1_state_0, TL04_jump_p1_state_1, TL04_jump_p2_state_0, TL04_jump_p2_state_1 : std_logic;
  signal TL04_n_0, TL04_n_1, TL04_n_2, TL04_n_4, TL04_n_5 : std_logic;
  signal TL04_n_6, TL04_n_7, TL04_n_8, TL04_n_9, TL04_n_10 : std_logic;
  signal TL04_n_11, TL04_n_12, TL04_n_13, TL04_n_14, TL04_n_15 : std_logic;
  signal TL04_n_16, TL04_n_17, TL04_n_18, TL04_n_19, TL04_n_20 : std_logic;
  signal TL04_n_21, TL04_n_22, TL04_n_23, TL04_n_24, TL04_n_25 : std_logic;
  signal TL04_n_26, TL04_n_27, TL04_n_28, TL04_n_29, TL04_n_30 : std_logic;
  signal TL04_n_31, TL04_n_33, TL04_n_36, TL04_n_37, TL04_n_38 : std_logic;
  signal UNCONNECTED, UNCONNECTED0, UNCONNECTED1, UNCONNECTED2, UNCONNECTED3 : std_logic;
  signal UNCONNECTED4, UNCONNECTED5, UNCONNECTED6, UNCONNECTED7, UNCONNECTED8 : std_logic;
  signal UNCONNECTED9, UNCONNECTED10, char1death, char2death, n_0 : std_logic;
  signal n_1, n_2, n_3, n_4, n_5 : std_logic;
  signal n_6, n_9, n_10, n_11, n_12 : std_logic;
  signal n_13, n_14, n_15, n_16, n_17 : std_logic;
  signal n_18, n_19, n_20, n_21, n_22 : std_logic;
  signal n_23, n_24, n_25, n_26, n_28 : std_logic;
  signal n_29, n_30, n_31, n_32, n_33 : std_logic;
  signal n_34, n_35, n_36, n_37, n_38 : std_logic;
  signal n_39, n_40, n_41, n_42, n_43 : std_logic;
  signal n_44, n_45, n_46, n_47, n_48 : std_logic;
  signal n_49, n_50, n_51, n_52, n_53 : std_logic;
  signal n_54, n_55, n_56, n_57, n_58 : std_logic;
  signal n_59, n_60, n_61, n_62, n_63 : std_logic;
  signal n_64, n_65, n_66, n_67, n_68 : std_logic;
  signal n_69, n_70, n_71, n_72, n_73 : std_logic;
  signal n_74, n_75, n_76, n_77, n_78 : std_logic;
  signal n_79, n_80, n_81, n_82, n_83 : std_logic;
  signal n_84, n_85, n_86, n_87, n_88 : std_logic;
  signal n_89, n_90, n_91, n_92, n_93 : std_logic;
  signal n_94, n_95, n_96, n_97, n_98 : std_logic;
  signal n_99, n_100, n_101, n_102, n_103 : std_logic;
  signal n_104, n_105, n_106, n_107, n_108 : std_logic;
  signal n_109, n_110, n_111, n_112, n_113 : std_logic;
  signal n_114, n_115, n_116, n_117, n_118 : std_logic;
  signal n_119, n_120, n_121, n_122, n_123 : std_logic;
  signal n_124, n_125, n_126, n_127, n_128 : std_logic;
  signal n_129, n_130, n_131, n_132, n_133 : std_logic;
  signal n_134, n_135, n_136, n_137, n_138 : std_logic;
  signal n_139, n_140, n_141, n_142, n_143 : std_logic;
  signal n_144, n_145, n_146, n_147, n_148 : std_logic;
  signal n_150, n_151, n_152, n_153, n_154 : std_logic;
  signal n_156, n_157, n_158, n_159, n_160 : std_logic;
  signal n_161, n_162, n_163, n_164, n_165 : std_logic;
  signal n_166, n_167, n_168, n_169, n_170 : std_logic;
  signal n_171, n_172, n_173, n_174, n_175 : std_logic;
  signal n_176, n_177, n_178, n_179, n_180 : std_logic;
  signal n_182, n_183, n_184, n_185, n_186 : std_logic;
  signal n_187, n_188, n_190, n_191, n_192 : std_logic;
  signal n_193, n_194, n_195, n_196, n_197 : std_logic;
  signal n_198, n_199, n_200, n_201, n_202 : std_logic;
  signal n_203, n_204, n_205, n_206, n_207 : std_logic;
  signal n_208, n_209, n_210, n_211, n_212 : std_logic;
  signal n_213, n_214, n_215, n_216, n_217 : std_logic;
  signal n_218, n_219, n_220, n_221, n_222 : std_logic;
  signal n_223, n_224, n_225, n_226, n_227 : std_logic;
  signal n_228, n_229, n_230, n_231, n_232 : std_logic;
  signal n_233, n_234, n_235, n_236, n_237 : std_logic;
  signal n_238, n_239, n_240, n_241, n_242 : std_logic;
  signal n_243, n_244, n_245, n_246, n_247 : std_logic;
  signal n_248, n_249, n_250, n_251, n_252 : std_logic;
  signal n_253, n_254, n_255, n_256, n_257 : std_logic;
  signal n_258, n_259, n_260, n_261, n_262 : std_logic;
  signal n_263, n_264, n_265, n_266, n_267 : std_logic;
  signal n_268, n_269, n_270, n_271, n_272 : std_logic;
  signal n_273, n_274, n_275, n_276, n_277 : std_logic;
  signal n_278, n_279, n_280, n_281, n_282 : std_logic;
  signal n_283, n_284, n_285, n_286, n_287 : std_logic;
  signal n_288, n_289, n_290, n_292, n_293 : std_logic;
  signal n_295, n_296, n_297, n_298, n_299 : std_logic;
  signal n_300, n_301, n_302, n_303, n_304 : std_logic;
  signal n_305, n_306, n_307, n_308, n_309 : std_logic;
  signal n_310, n_311, n_312, n_313, n_314 : std_logic;
  signal n_315, n_316, n_317, n_318, n_319 : std_logic;
  signal n_320, n_321, n_322, n_323, n_324 : std_logic;
  signal n_325, n_326, n_327, n_328, n_329 : std_logic;
  signal n_330, n_331, n_332, n_333, n_334 : std_logic;
  signal n_335, n_336, n_337, n_338, n_339 : std_logic;
  signal n_340, n_341, n_342, n_343, n_344 : std_logic;
  signal n_345, n_346, n_347, n_348, n_349 : std_logic;
  signal n_350, n_351, n_352, n_353, n_354 : std_logic;
  signal n_355, n_356, n_357, n_358, n_359 : std_logic;
  signal n_360, n_361, n_362, n_363, n_364 : std_logic;
  signal n_365, n_366, n_367, n_368, n_369 : std_logic;
  signal n_370, n_371, n_372, n_373, n_374 : std_logic;
  signal n_375, n_376, n_377, n_378, n_379 : std_logic;
  signal n_380, n_381, n_382, n_383, n_384 : std_logic;
  signal n_385, n_386, n_387, n_389, n_390 : std_logic;
  signal n_391, n_392, n_393, n_395, n_396 : std_logic;
  signal n_397, n_398, n_399, n_400, n_401 : std_logic;
  signal n_402, n_403, n_404, n_405, n_406 : std_logic;
  signal n_407, n_408, n_409, n_410, n_411 : std_logic;
  signal n_412, n_413, n_414, n_415, n_416 : std_logic;
  signal n_417, n_418, n_419, n_420, n_421 : std_logic;
  signal n_422, n_423, n_424, n_425, n_426 : std_logic;
  signal n_427, n_428, n_429, n_430, n_431 : std_logic;
  signal n_432, n_433, n_434, n_435, n_436 : std_logic;
  signal n_437, n_438, n_439, n_440, n_441 : std_logic;
  signal n_442, n_443, n_444, n_445, n_446 : std_logic;
  signal n_447, n_448, n_449, n_450, n_451 : std_logic;
  signal n_452, n_453, n_454, n_455, n_456 : std_logic;
  signal n_457, n_458, n_459, n_460, n_461 : std_logic;
  signal n_462, n_463, n_464, n_465, n_466 : std_logic;
  signal n_467, n_468, n_469, n_470, n_471 : std_logic;
  signal n_472, n_473, n_474, n_478, n_479 : std_logic;
  signal n_480, n_482, n_483, n_484, n_485 : std_logic;
  signal n_487, n_504, n_505, n_506, n_507 : std_logic;
  signal n_508, orientationp1, orientationp2 : std_logic;

begin

  B_data(2) <= G_data(3);
  G_data(1) <= R_data(1);
  R_data(2) <= R_data(3);
  FE_PHC177_char1posyin_1 : DEL01BWP7T port map(I => FE_PHN159_char1posyin_1, Z => FE_PHN177_char1posyin_1);
  FE_PHC176_char2velx_9 : DEL01BWP7T port map(I => char2velx(9), Z => FE_PHN176_char2velx_9);
  FE_PHC175_char2vely_3 : DEL01BWP7T port map(I => FE_PHN175_char2vely_3, Z => char2vely(3));
  FE_PHC174_vcountintern_8 : DEL01BWP7T port map(I => vcountintern(8), Z => FE_PHN174_vcountintern_8);
  FE_PHC173_TL04_driver_pulse_count_0 : DEL01BWP7T port map(I => TL04_driver_pulse_count_0, Z => FE_PHN173_TL04_driver_pulse_count_0);
  FE_PHC172_TL01_CLR1_n_1491 : DEL01BWP7T port map(I => TL01_CLR1_n_1491, Z => FE_PHN172_TL01_CLR1_n_1491);
  FE_PHC171_TL01_CLR1_char2_sprite_frame_control_frame_count_2 : DEL01BWP7T port map(I => TL01_CLR1_char2_sprite_frame_control_frame_count_2, Z => FE_PHN171_TL01_CLR1_char2_sprite_frame_control_frame_count_2);
  FE_PHC170_TL04_n_15 : DEL01BWP7T port map(I => FE_PHN155_TL04_n_15, Z => FE_PHN170_TL04_n_15);
  FE_PHC169_TL01_CLR1_char2_sprite_frame_control_cnt_reset : CKBD0BWP7T port map(I => FE_PHN60_TL01_CLR1_char2_sprite_frame_control_cnt_reset, Z => FE_PHN169_TL01_CLR1_char2_sprite_frame_control_cnt_reset);
  FE_PHC168_char2posy_7 : DEL01BWP7T port map(I => FE_PHN91_char2posy_7, Z => FE_PHN168_char2posy_7);
  FE_PHC167_char1posxin_5 : DEL01BWP7T port map(I => FE_PHN69_char1posxin_5, Z => FE_PHN167_char1posxin_5);
  FE_PHC166_TL01_CLR1_char1_sprite_frame_control_cnt_reset : DEL01BWP7T port map(I => TL01_CLR1_char1_sprite_frame_control_cnt_reset, Z => FE_PHN166_TL01_CLR1_char1_sprite_frame_control_cnt_reset);
  FE_PHC165_char2posx_1 : DEL01BWP7T port map(I => FE_PHN94_char2posx_1, Z => FE_PHN165_char2posx_1);
  FE_PHC164_char2posx_0 : DEL01BWP7T port map(I => FE_PHN92_char2posx_0, Z => FE_PHN164_char2posx_0);
  FE_PHC163_TL01_CLR1_char2_sprite_frame_control_frame_count_4 : DEL01BWP7T port map(I => TL01_CLR1_char2_sprite_frame_control_frame_count_4, Z => FE_PHN163_TL01_CLR1_char2_sprite_frame_control_frame_count_4);
  FE_PHC162_char1posxin_6 : DEL01BWP7T port map(I => FE_PHN67_char1posxin_6, Z => FE_PHN162_char1posxin_6);
  FE_PHC161_TL01_CLR1_char1_sprite_frame_control_frame_count_0 : DEL01BWP7T port map(I => TL01_CLR1_char1_sprite_frame_control_frame_count_0, Z => FE_PHN161_TL01_CLR1_char1_sprite_frame_control_frame_count_0);
  FE_PHC160_TL01_SCNR1_hcount_reset : DEL01BWP7T port map(I => FE_PHN68_TL01_SCNR1_hcount_reset, Z => FE_PHN160_TL01_SCNR1_hcount_reset);
  FE_PHC159_char1posyin_1 : CKBD0BWP7T port map(I => char1posyin(1), Z => FE_PHN159_char1posyin_1);
  FE_PHC158_TL01_n_0 : DEL01BWP7T port map(I => TL01_n_0, Z => FE_PHN158_TL01_n_0);
  FE_PHC157_ATT1_n_34 : DEL1BWP7T port map(I => ATT1_n_34, Z => FE_PHN157_ATT1_n_34);
  FE_PHC156_ATT1_n_26 : DEL0BWP7T port map(I => ATT1_n_26, Z => FE_PHN156_ATT1_n_26);
  FE_PHC155_TL04_n_15 : CKBD0BWP7T port map(I => TL04_n_15, Z => FE_PHN155_TL04_n_15);
  FE_PHC154_TL01_CLR1_n_33 : CKBD0BWP7T port map(I => TL01_CLR1_n_33, Z => FE_PHN154_TL01_CLR1_n_33);
  FE_PHC153_TL01_CLR1_n_41 : CKBD0BWP7T port map(I => TL01_CLR1_n_41, Z => FE_PHN153_TL01_CLR1_n_41);
  FE_PHC152_TL01_CLR1_n_303 : DEL02BWP7T port map(I => TL01_CLR1_n_303, Z => FE_PHN152_TL01_CLR1_n_303);
  FE_PHC151_TL01_CLR1_n_32 : DEL0BWP7T port map(I => FE_PHN151_TL01_CLR1_n_32, Z => TL01_CLR1_n_32);
  FE_PHC150_TL01_CLR1_n_34 : DEL0BWP7T port map(I => TL01_CLR1_n_34, Z => FE_PHN150_TL01_CLR1_n_34);
  FE_PHC149_TL01_CLR1_n_305 : DEL0BWP7T port map(I => FE_PHN149_TL01_CLR1_n_305, Z => TL01_CLR1_n_305);
  FE_PHC148_ATT1_n_32 : DEL1BWP7T port map(I => FE_PHN148_ATT1_n_32, Z => ATT1_n_32);
  FE_PHC147_TL01_CLR1_n_257 : DEL01BWP7T port map(I => TL01_CLR1_n_257, Z => FE_PHN147_TL01_CLR1_n_257);
  FE_PHC146_ATT1_n_12 : DEL0BWP7T port map(I => ATT1_n_12, Z => FE_PHN146_ATT1_n_12);
  FE_PHC145_ATT1_n_35 : DEL0BWP7T port map(I => ATT1_n_35, Z => FE_PHN145_ATT1_n_35);
  FE_PHC144_TL01_CLR1_n_733 : DEL0BWP7T port map(I => TL01_CLR1_n_733, Z => FE_PHN144_TL01_CLR1_n_733);
  FE_PHC143_n_73 : DEL0BWP7T port map(I => FE_PHN143_n_73, Z => n_73);
  FE_PHC142_n_108 : DEL0BWP7T port map(I => n_108, Z => FE_PHN142_n_108);
  FE_PHC141_n_109 : DEL0BWP7T port map(I => n_109, Z => FE_PHN141_n_109);
  FE_PHC140_n_101 : DEL0BWP7T port map(I => FE_PHN140_n_101, Z => n_101);
  FE_PHC139_n_74 : DEL0BWP7T port map(I => n_74, Z => FE_PHN139_n_74);
  FE_PHC138_n_71 : DEL0BWP7T port map(I => FE_PHN138_n_71, Z => n_71);
  FE_PHC137_n_111 : DEL0BWP7T port map(I => n_111, Z => FE_PHN137_n_111);
  FE_PHC136_n_107 : DEL0BWP7T port map(I => FE_PHN136_n_107, Z => n_107);
  FE_PHC135_n_99 : DEL0BWP7T port map(I => n_99, Z => FE_PHN135_n_99);
  FE_PHC134_n_72 : DEL0BWP7T port map(I => n_72, Z => FE_PHN134_n_72);
  FE_PHC133_n_70 : DEL0BWP7T port map(I => n_70, Z => FE_PHN133_n_70);
  FE_PHC132_n_75 : DEL0BWP7T port map(I => n_75, Z => FE_PHN132_n_75);
  FE_PHC131_n_105 : DEL0BWP7T port map(I => n_105, Z => FE_PHN131_n_105);
  FE_PHC130_n_98 : DEL0BWP7T port map(I => n_98, Z => FE_PHN130_n_98);
  FE_PHC129_TL04_n_23 : DEL0BWP7T port map(I => FE_PHN129_TL04_n_23, Z => TL04_n_23);
  FE_PHC128_n_113 : DEL0BWP7T port map(I => n_113, Z => FE_PHN128_n_113);
  FE_PHC127_n_88 : DEL0BWP7T port map(I => n_88, Z => FE_PHN127_n_88);
  FE_PHC126_ATT1_n_25 : DEL0BWP7T port map(I => ATT1_n_25, Z => FE_PHN126_ATT1_n_25);
  FE_PHC125_TL04_n_27 : DEL0BWP7T port map(I => TL04_n_27, Z => FE_PHN125_TL04_n_27);
  FE_PHC124_char1posx_8 : CKBD0BWP7T port map(I => FE_PHN124_char1posx_8, Z => char1posx(8));
  FE_PHC123_char2posx_8 : CKBD0BWP7T port map(I => char2posx(8), Z => FE_PHN123_char2posx_8);
  FE_PHC122_vcountintern_9 : CKBD0BWP7T port map(I => FE_PHN122_vcountintern_9, Z => vcountintern(9));
  FE_PHC121_ATT1_PM2_state2_1 : DEL02BWP7T port map(I => FE_PHN121_ATT1_PM2_state2_1, Z => ATT1_PM2_state2_1);
  FE_PHC120_ATT1_PM2_state2_0 : DEL02BWP7T port map(I => FE_PHN120_ATT1_PM2_state2_0, Z => ATT1_PM2_state2_0);
  FE_PHC119_char2posx_6 : DEL01BWP7T port map(I => char2posx(6), Z => FE_PHN119_char2posx_6);
  FE_PHC118_char2perc_1 : DEL01BWP7T port map(I => char2perc(1), Z => FE_PHN118_char2perc_1);
  FE_PHC117_char2perc_7 : DEL01BWP7T port map(I => char2perc(7), Z => FE_PHN117_char2perc_7);
  FE_PHC116_ATT1_PM2_state1_1 : DEL02BWP7T port map(I => ATT1_PM2_state1_1, Z => FE_PHN116_ATT1_PM2_state1_1);
  FE_PHC115_ATT1_PM4_state2_1 : DEL0BWP7T port map(I => FE_PHN115_ATT1_PM4_state2_1, Z => ATT1_PM4_state2_1);
  FE_PHC114_ATT1_PM4_state2_0 : DEL0BWP7T port map(I => FE_PHN114_ATT1_PM4_state2_0, Z => ATT1_PM4_state2_0);
  FE_PHC113_TL04_driver_state_0 : DEL02BWP7T port map(I => TL04_driver_state_0, Z => FE_PHN113_TL04_driver_state_0);
  FE_PHC112_char1perc_7 : DEL01BWP7T port map(I => char1perc(7), Z => FE_PHN112_char1perc_7);
  FE_PHC111_TL01_CLR1_char1_sprite_frame_control_frame_count_2 : CKBD0BWP7T port map(I => TL01_CLR1_char1_sprite_frame_control_frame_count_2, Z => FE_PHN111_TL01_CLR1_char1_sprite_frame_control_frame_count_2);
  FE_PHC110_char1perc_0 : DEL01BWP7T port map(I => char1perc(0), Z => FE_PHN110_char1perc_0);
  FE_PHC109_TL01_CLR1_char1_sprite_frame_control_frame_count_3 : DEL02BWP7T port map(I => TL01_CLR1_char1_sprite_frame_control_frame_count_3, Z => FE_PHN109_TL01_CLR1_char1_sprite_frame_control_frame_count_3);
  FE_PHC108_TL01_CLR1_char1_sprite_frame_control_frame_count_0 : DEL02BWP7T port map(I => FE_PHN108_TL01_CLR1_char1_sprite_frame_control_frame_count_0, Z => TL01_CLR1_char1_sprite_frame_control_frame_count_0);
  FE_PHC107_TL01_CLR1_char2_sprite_frame_control_frame_count_0 : DEL0BWP7T port map(I => FE_PHN107_TL01_CLR1_char2_sprite_frame_control_frame_count_0, Z => TL01_CLR1_char2_sprite_frame_control_frame_count_0);
  FE_PHC106_TL01_CLR1_char1_sprite_frame_control_state_0 : CKBD0BWP7T port map(I => TL01_CLR1_char1_sprite_frame_control_state_0, Z => FE_PHN106_TL01_CLR1_char1_sprite_frame_control_state_0);
  FE_PHC105_TL01_CLR1_char1_sprite_frame_control_frame_count_4 : DEL02BWP7T port map(I => FE_PHN105_TL01_CLR1_char1_sprite_frame_control_frame_count_4, Z => TL01_CLR1_char1_sprite_frame_control_frame_count_4);
  FE_PHC104_TL04_driver_state_1 : CKBD0BWP7T port map(I => FE_PHN104_TL04_driver_state_1, Z => TL04_driver_state_1);
  FE_PHC103_TL01_CLR1_char1_sprite_frame_control_state_2 : CKBD0BWP7T port map(I => FE_PHN103_TL01_CLR1_char1_sprite_frame_control_state_2, Z => TL01_CLR1_char1_sprite_frame_control_state_2);
  FE_PHC102_char2perc_0 : DEL01BWP7T port map(I => char2perc(0), Z => FE_PHN102_char2perc_0);
  FE_PHC101_char2posy_2 : DEL01BWP7T port map(I => char2posy(2), Z => FE_PHN101_char2posy_2);
  FE_PHC100_char2posx_3 : DEL01BWP7T port map(I => char2posx(3), Z => FE_PHN100_char2posx_3);
  FE_PHC99_TL01_CLR1_char2_sprite_frame_control_state_2 : CKBD0BWP7T port map(I => TL01_CLR1_char2_sprite_frame_control_state_2, Z => FE_PHN99_TL01_CLR1_char2_sprite_frame_control_state_2);
  FE_PHC98_inputsp2_5 : DEL0BWP7T port map(I => inputsp2(5), Z => FE_PHN98_inputsp2_5);
  FE_PHC97_char2perc_2 : CKBD0BWP7T port map(I => char2perc(2), Z => FE_PHN97_char2perc_2);
  FE_PHC96_TL01_n_1 : DEL01BWP7T port map(I => TL01_n_1, Z => FE_PHN96_TL01_n_1);
  FE_PHC95_char2posy_0 : DEL0BWP7T port map(I => char2posy(0), Z => FE_PHN95_char2posy_0);
  FE_PHC94_char2posx_1 : CKBD0BWP7T port map(I => char2posx(1), Z => FE_PHN94_char2posx_1);
  FE_PHC93_char2posy_6 : DEL01BWP7T port map(I => char2posy(6), Z => FE_PHN93_char2posy_6);
  FE_PHC92_char2posx_0 : CKBD0BWP7T port map(I => char2posx(0), Z => FE_PHN92_char2posx_0);
  FE_PHC91_char2posy_7 : CKBD0BWP7T port map(I => char2posy(7), Z => FE_PHN91_char2posy_7);
  FE_PHC90_char2perc_3 : CKBD0BWP7T port map(I => char2perc(3), Z => FE_PHN90_char2perc_3);
  FE_PHC89_TL04_n_0 : DEL01BWP7T port map(I => TL04_n_0, Z => FE_PHN89_TL04_n_0);
  FE_PHC88_TL01_CLR1_char2_sprite_frame_control_state_0 : DEL02BWP7T port map(I => FE_PHN88_TL01_CLR1_char2_sprite_frame_control_state_0, Z => TL01_CLR1_char2_sprite_frame_control_state_0);
  FE_PHC87_char2velx_9 : CKBD0BWP7T port map(I => FE_PHN176_char2velx_9, Z => FE_PHN87_char2velx_9);
  FE_PHC86_char2vely_3 : CKBD0BWP7T port map(I => char2vely(3), Z => FE_PHN86_char2vely_3);
  FE_PHC85_char2posx_2 : CKBD0BWP7T port map(I => char2posx(2), Z => FE_PHN85_char2posx_2);
  FE_PHC84_TL01_CLR1_char2_sprite_frame_control_frame_count_3 : DEL02BWP7T port map(I => TL01_CLR1_char2_sprite_frame_control_frame_count_3, Z => FE_PHN84_TL01_CLR1_char2_sprite_frame_control_frame_count_3);
  FE_PHC83_char2posy_3 : DEL0BWP7T port map(I => char2posy(3), Z => FE_PHN83_char2posy_3);
  FE_PHC82_char2posx_4 : CKBD0BWP7T port map(I => char2posx(4), Z => FE_PHN82_char2posx_4);
  FE_PHC81_char2posy_1 : DEL0BWP7T port map(I => char2posy(1), Z => FE_PHN81_char2posy_1);
  FE_PHC80_TL04_driver_pulse_count_0 : DEL02BWP7T port map(I => FE_PHN80_TL04_driver_pulse_count_0, Z => TL04_driver_pulse_count_0);
  FE_PHC79_char2posy_4 : CKBD0BWP7T port map(I => char2posy(4), Z => FE_PHN79_char2posy_4);
  FE_PHC78_TL04_n_11 : DEL0BWP7T port map(I => TL04_n_11, Z => FE_PHN78_TL04_n_11);
  FE_PHC77_char2velx_1 : DEL0BWP7T port map(I => char2velx(1), Z => FE_PHN77_char2velx_1);
  FE_PHC76_char2velx_3 : DEL0BWP7T port map(I => char2velx(3), Z => FE_PHN76_char2velx_3);
  FE_PHC75_char2velx_4 : DEL0BWP7T port map(I => char2velx(4), Z => FE_PHN75_char2velx_4);
  FE_PHC74_TL04_n_13 : DEL0BWP7T port map(I => TL04_n_13, Z => FE_PHN74_TL04_n_13);
  FE_PHC73_char2velx_0 : DEL0BWP7T port map(I => char2velx(0), Z => FE_PHN73_char2velx_0);
  FE_PHC72_char2posy_5 : CKBD0BWP7T port map(I => char2posy(5), Z => FE_PHN72_char2posy_5);
  FE_PHC71_char2velx_2 : DEL0BWP7T port map(I => char2velx(2), Z => FE_PHN71_char2velx_2);
  FE_PHC70_char2velx_7 : DEL0BWP7T port map(I => char2velx(7), Z => FE_PHN70_char2velx_7);
  FE_PHC69_char1posxin_5 : DEL02BWP7T port map(I => char1posxin(5), Z => FE_PHN69_char1posxin_5);
  FE_PHC68_TL01_SCNR1_hcount_reset : CKBD0BWP7T port map(I => TL01_SCNR1_hcount_reset, Z => FE_PHN68_TL01_SCNR1_hcount_reset);
  FE_PHC67_char1posxin_6 : DEL02BWP7T port map(I => char1posxin(6), Z => FE_PHN67_char1posxin_6);
  FE_PHC66_char2velx_5 : DEL0BWP7T port map(I => char2velx(5), Z => FE_PHN66_char2velx_5);
  FE_PHC65_TL04_n_10 : DEL0BWP7T port map(I => TL04_n_10, Z => FE_PHN65_TL04_n_10);
  FE_PHC64_TL04_n_12 : DEL0BWP7T port map(I => TL04_n_12, Z => FE_PHN64_TL04_n_12);
  FE_PHC63_char1posyin_1 : DEL02BWP7T port map(I => FE_PHN63_char1posyin_1, Z => char1posyin(1));
  FE_PHC62_TL01_n_0 : DEL02BWP7T port map(I => FE_PHN62_TL01_n_0, Z => TL01_n_0);
  FE_PHC61_char1velxin_8 : DEL2BWP7T port map(I => char1velxin(8), Z => FE_PHN61_char1velxin_8);
  FE_PHC60_TL01_CLR1_char2_sprite_frame_control_cnt_reset : DEL02BWP7T port map(I => TL01_CLR1_char2_sprite_frame_control_cnt_reset, Z => FE_PHN60_TL01_CLR1_char2_sprite_frame_control_cnt_reset);
  FE_PHC59_TL01_CLR1_char1_sprite_frame_control_cnt_reset : DEL02BWP7T port map(I => FE_PHN166_TL01_CLR1_char1_sprite_frame_control_cnt_reset, Z => FE_PHN59_TL01_CLR1_char1_sprite_frame_control_cnt_reset);
  FE_PHC58_TL00_WL00_state_1 : DEL2BWP7T port map(I => TL00_WL00_state_1, Z => FE_PHN58_TL00_WL00_state_1);
  FE_PHC57_char1posxin_7 : DEL0BWP7T port map(I => FE_PHN57_char1posxin_7, Z => char1posxin(7));
  FE_PHC56_char1posxin_2 : DEL0BWP7T port map(I => FE_PHN56_char1posxin_2, Z => char1posxin(2));
  FE_PHC55_char1posxin_1 : DEL0BWP7T port map(I => char1posxin(1), Z => FE_PHN55_char1posxin_1);
  FE_PHC54_char1posxin_3 : DEL0BWP7T port map(I => char1posxin(3), Z => FE_PHN54_char1posxin_3);
  FE_PHC53_TL01_CLR1_n_1 : DEL0BWP7T port map(I => TL01_CLR1_n_1, Z => FE_PHN53_TL01_CLR1_n_1);
  FE_PHC52_char1posxin_8 : DEL0BWP7T port map(I => char1posxin(8), Z => FE_PHN52_char1posxin_8);
  FE_PHC51_TL01_CLR1_n_0 : DEL0BWP7T port map(I => FE_PHN51_TL01_CLR1_n_0, Z => TL01_CLR1_n_0);
  FE_PHC50_char1posxin_4 : DEL0BWP7T port map(I => char1posxin(4), Z => FE_PHN50_char1posxin_4);
  FE_PHC49_char1posxin_0 : DEL0BWP7T port map(I => FE_PHN49_char1posxin_0, Z => char1posxin(0));
  FE_PHC48_ATT1_n_5 : DEL0BWP7T port map(I => FE_PHN48_ATT1_n_5, Z => ATT1_n_5);
  FE_PHC47_char1posyin_2 : DEL0BWP7T port map(I => FE_PHN47_char1posyin_2, Z => char1posyin(2));
  FE_PHC46_char1posyin_7 : DEL0BWP7T port map(I => char1posyin(7), Z => FE_PHN46_char1posyin_7);
  FE_PHC45_char1posyin_6 : DEL0BWP7T port map(I => FE_PHN45_char1posyin_6, Z => char1posyin(6));
  FE_PHC44_char1posyin_3 : DEL0BWP7T port map(I => FE_PHN44_char1posyin_3, Z => char1posyin(3));
  FE_PHC43_char1posyin_5 : DEL0BWP7T port map(I => FE_PHN43_char1posyin_5, Z => char1posyin(5));
  FE_PHC42_char1posyin_4 : DEL0BWP7T port map(I => FE_PHN42_char1posyin_4, Z => char1posyin(4));
  FE_PHC41_char1posyin_0 : DEL0BWP7T port map(I => FE_PHN41_char1posyin_0, Z => char1posyin(0));
  FE_PHC40_char1velyin_9 : DEL0BWP7T port map(I => FE_PHN40_char1velyin_9, Z => char1velyin(9));
  FE_PHC39_char1velyin_6 : DEL0BWP7T port map(I => char1velyin(6), Z => FE_PHN39_char1velyin_6);
  FE_PHC38_char1velyin_8 : DEL0BWP7T port map(I => FE_PHN38_char1velyin_8, Z => char1velyin(8));
  FE_PHC37_char1velyin_7 : DEL0BWP7T port map(I => FE_PHN37_char1velyin_7, Z => char1velyin(7));
  FE_PHC36_char1velxin_6 : DEL0BWP7T port map(I => FE_PHN36_char1velxin_6, Z => char1velxin(6));
  FE_PHC35_char1velyin_1 : DEL0BWP7T port map(I => FE_PHN35_char1velyin_1, Z => char1velyin(1));
  FE_PHC34_TL01_n_2 : CKBD0BWP7T port map(I => FE_PHN34_TL01_n_2, Z => TL01_n_2);
  FE_PHC33_char1velyin_0 : DEL0BWP7T port map(I => FE_PHN33_char1velyin_0, Z => char1velyin(0));
  FE_PHC32_char1velxin_0 : DEL0BWP7T port map(I => char1velxin(0), Z => FE_PHN32_char1velxin_0);
  FE_PHC31_char1velyin_4 : DEL0BWP7T port map(I => char1velyin(4), Z => FE_PHN31_char1velyin_4);
  FE_PHC30_char1velyin_2 : DEL0BWP7T port map(I => char1velyin(2), Z => FE_PHN30_char1velyin_2);
  FE_PHC29_char1velxin_1 : DEL0BWP7T port map(I => FE_PHN29_char1velxin_1, Z => char1velxin(1));
  FE_PHC28_char1velyin_5 : DEL0BWP7T port map(I => FE_PHN28_char1velyin_5, Z => char1velyin(5));
  FE_PHC27_char1velxin_5 : DEL0BWP7T port map(I => char1velxin(5), Z => FE_PHN27_char1velxin_5);
  FE_PHC26_char1velxin_3 : DEL0BWP7T port map(I => FE_PHN26_char1velxin_3, Z => char1velxin(3));
  FE_PHC25_char1velxin_2 : DEL0BWP7T port map(I => char1velxin(2), Z => FE_PHN25_char1velxin_2);
  FE_PHC24_char1velyin_3 : DEL0BWP7T port map(I => char1velyin(3), Z => FE_PHN24_char1velyin_3);
  FE_PHC23_char1velxin_7 : DEL0BWP7T port map(I => FE_PHN23_char1velxin_7, Z => char1velxin(7));
  FE_PHC22_char1velxin_4 : DEL0BWP7T port map(I => char1velxin(4), Z => FE_PHN22_char1velxin_4);
  FE_PHC21_char1velxin_9 : DEL0BWP7T port map(I => char1velxin(9), Z => FE_PHN21_char1velxin_9);
  FE_PHC20_TL01_CLR1_char2_sprite_frame_control_new_state_0 : DEL1BWP7T port map(I => TL01_CLR1_char2_sprite_frame_control_new_state_0, Z => FE_PHN20_TL01_CLR1_char2_sprite_frame_control_new_state_0);
  FE_PHC19_TL01_CLR1_char1_sprite_frame_control_new_state_0 : DEL1BWP7T port map(I => TL01_CLR1_char1_sprite_frame_control_new_state_0, Z => FE_PHN19_TL01_CLR1_char1_sprite_frame_control_new_state_0);
  FE_PHC18_TL01_CLR1_char2_sprite_frame_control_new_state_1 : DEL1BWP7T port map(I => TL01_CLR1_char2_sprite_frame_control_new_state_1, Z => FE_PHN18_TL01_CLR1_char2_sprite_frame_control_new_state_1);
  FE_PHC17_TL01_CLR1_char2_sprite_frame_control_new_state_2 : DEL1BWP7T port map(I => TL01_CLR1_char2_sprite_frame_control_new_state_2, Z => FE_PHN17_TL01_CLR1_char2_sprite_frame_control_new_state_2);
  FE_PHC16_TL01_CLR1_char1_sprite_frame_control_new_state_1 : DEL1BWP7T port map(I => TL01_CLR1_char1_sprite_frame_control_new_state_1, Z => FE_PHN16_TL01_CLR1_char1_sprite_frame_control_new_state_1);
  FE_PHC15_TL01_CLR1_char1_sprite_frame_control_new_state_2 : DEL1BWP7T port map(I => TL01_CLR1_char1_sprite_frame_control_new_state_2, Z => FE_PHN15_TL01_CLR1_char1_sprite_frame_control_new_state_2);
  FE_OFC4_TL00_writeint : BUFFD1P5BWP7T port map(I => TL00_writeint, Z => FE_OFN4_TL00_writeint);
  FE_OFC3_reset : DEL01BWP7T port map(I => reset, Z => FE_OFN3_reset);
  FE_OFC2_ATT1_n_301 : DEL01BWP7T port map(I => ATT1_n_301, Z => FE_OFN2_ATT1_n_301);
  FE_OFC1_TL02_PHS0_sel_0 : BUFFD2BWP7T port map(I => TL02_PHS0_sel_0, Z => FE_OFN1_TL02_PHS0_sel_0);
  FE_OFC0_n_6 : BUFFD2BWP7T port map(I => n_6, Z => FE_OFN0_n_6);
  CTS_ccl_a_BUF_clk_G0_L2_3 : CKBD12BWP7T port map(I => CTS_18, Z => CTS_17);
  CTS_ccl_a_BUF_clk_G0_L2_2 : CKBD12BWP7T port map(I => CTS_18, Z => CTS_16);
  CTS_ccl_a_BUF_clk_G0_L2_1 : CKBD12BWP7T port map(I => CTS_18, Z => CTS_15);
  CTS_ccl_a_BUF_clk_G0_L1_1 : CKBD8BWP7T port map(I => clk, Z => CTS_18);
  FE_DBTC14_reset : INVD2BWP7T port map(I => FE_OFN3_reset, ZN => FE_DBTN14_reset);
  FE_DBTC13_char1perc_5 : INVD1BWP7T port map(I => char1perc(5), ZN => FE_DBTN13_char1perc_5);
  FE_DBTC12_char1perc_4 : INVD1BWP7T port map(I => char1perc(4), ZN => FE_DBTN12_char1perc_4);
  FE_DBTC11_char1perc_3 : INVD0BWP7T port map(I => char1perc(3), ZN => FE_DBTN11_char1perc_3);
  FE_DBTC10_char1perc_1 : INVD0BWP7T port map(I => char1perc(1), ZN => FE_DBTN10_char1perc_1);
  FE_DBTC9_char2perc_5 : INVD1BWP7T port map(I => char2perc(5), ZN => FE_DBTN9_char2perc_5);
  FE_DBTC8_char2perc_4 : INVD1BWP7T port map(I => char2perc(4), ZN => FE_DBTN8_char2perc_4);
  FE_DBTC7_char2perc_3 : INVD1BWP7T port map(I => char2perc(3), ZN => FE_DBTN7_char2perc_3);
  FE_DBTC6_char2perc_2 : INVD1BWP7T port map(I => char2perc(2), ZN => FE_DBTN6_char2perc_2);
  FE_DBTC5_char2perc_1 : INVD1BWP7T port map(I => char2perc(1), ZN => FE_DBTN5_char2perc_1);
  FE_DBTC4_char2perc_0 : INVD0BWP7T port map(I => char2perc(0), ZN => FE_DBTN4_char2perc_0);
  FE_DBTC3_char1posx_4 : INVD0BWP7T port map(I => char1posx(4), ZN => FE_DBTN3_char1posx_4);
  FE_DBTC2_char1posy_3 : INVD1BWP7T port map(I => char1posy(3), ZN => FE_DBTN2_char1posy_3);
  FE_DBTC1_char2posx_1 : INVD0BWP7T port map(I => char2posx(1), ZN => FE_DBTN1_char2posx_1);
  FE_DBTC0_char2posx_0 : INVD0BWP7T port map(I => char2posx(0), ZN => FE_DBTN0_char2posx_0);
  ATT1_PM1 : orientation port map(clk => clk, res => reset, input1 => inputsp1, input2 => inputsp2, output1 => orientationp1, output2 => orientationp2);
  TL04_counter : input_period_counter port map(clk => clk, reset => TL04_count_reset, count_out => TL04_count);
  g646 : IAO21D0BWP7T port map(A1 => n_485, A2 => TL02_kb_y_5, B => TL02_kb_y_6, ZN => n_487);
  g647 : OR4D1BWP7T port map(A1 => TL02_kb_y_4, A2 => TL02_kb_y_3, A3 => TL02_kb_y_1, A4 => n_484, Z => n_485);
  g648 : IND3D1BWP7T port map(A1 => TL02_kb_y_2, B1 => n_482, B2 => n_483, ZN => n_484);
  g649 : INVD1BWP7T port map(I => n_483, ZN => TL02_kb_y_0);
  g650 : AO22D0BWP7T port map(A1 => FE_OFN1_TL02_PHS0_sel_0, A2 => dirx2new2(1), B1 => FE_OFN0_n_6, B2 => dirx1new2(1), Z => TL02_n_444);
  g651 : AO22D0BWP7T port map(A1 => char1perctemp(6), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => char2perctemp(6), Z => TL02_n_447);
  g652 : AO22D0BWP7T port map(A1 => FE_OFN0_n_6, A2 => dirx1new2(4), B1 => dirx2new2(4), B2 => FE_OFN1_TL02_PHS0_sel_0, Z => TL02_n_441);
  g653 : AO22D0BWP7T port map(A1 => FE_OFN0_n_6, A2 => dirx1new2(3), B1 => dirx2new2(3), B2 => FE_OFN1_TL02_PHS0_sel_0, Z => TL02_n_442);
  g654 : AO22D0BWP7T port map(A1 => FE_OFN0_n_6, A2 => dirx1new2(2), B1 => dirx2new2(2), B2 => FE_OFN1_TL02_PHS0_sel_0, Z => TL02_n_443);
  g655 : AO22D0BWP7T port map(A1 => char1perctemp(7), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => char2perctemp(7), Z => TL02_n_446);
  g656 : AOI22D0BWP7T port map(A1 => FE_OFN0_n_6, A2 => diry1new2(7), B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => diry2new2(7), ZN => n_482);
  g657 : AO22D0BWP7T port map(A1 => dirx1new2(0), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => dirx2new2(0), Z => TL02_n_445);
  g658 : AO22D0BWP7T port map(A1 => diry1new2(2), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => diry2new2(2), Z => TL02_kb_y_2);
  g659 : AO22D0BWP7T port map(A1 => FE_OFN1_TL02_PHS0_sel_0, A2 => diry2new2(5), B1 => FE_OFN0_n_6, B2 => diry1new2(5), Z => TL02_kb_y_5);
  g660 : AO22D0BWP7T port map(A1 => diry1new2(3), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => diry2new2(3), Z => TL02_kb_y_3);
  g661 : AOI22D0BWP7T port map(A1 => diry1new2(0), A2 => FE_OFN0_n_6, B1 => diry2new2(0), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_483);
  g662 : AO22D0BWP7T port map(A1 => char1perctemp(0), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => char2perctemp(0), Z => TL02_n_453);
  g663 : AO22D0BWP7T port map(A1 => char1perctemp(4), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => char2perctemp(4), Z => TL02_n_449);
  g664 : AO22D0BWP7T port map(A1 => FE_OFN0_n_6, A2 => dirx1new2(6), B1 => dirx2new2(6), B2 => FE_OFN1_TL02_PHS0_sel_0, Z => TL02_n_439);
  g665 : AO22D0BWP7T port map(A1 => char1perctemp(3), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => char2perctemp(3), Z => TL02_n_450);
  g666 : AO22D0BWP7T port map(A1 => FE_OFN0_n_6, A2 => dirx1new2(7), B1 => dirx2new2(7), B2 => FE_OFN1_TL02_PHS0_sel_0, Z => TL02_n_438);
  g667 : AO22D0BWP7T port map(A1 => FE_OFN0_n_6, A2 => dirx1new2(5), B1 => dirx2new2(5), B2 => FE_OFN1_TL02_PHS0_sel_0, Z => TL02_n_440);
  g668 : AO22D0BWP7T port map(A1 => char1perctemp(2), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => char2perctemp(2), Z => TL02_n_451);
  g669 : AO22D0BWP7T port map(A1 => char1perctemp(1), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => char2perctemp(1), Z => TL02_n_452);
  g670 : AO22D0BWP7T port map(A1 => char1perctemp(5), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => char2perctemp(5), Z => TL02_n_448);
  g671 : AO22D0BWP7T port map(A1 => FE_OFN0_n_6, A2 => diry1new2(6), B1 => diry2new2(6), B2 => FE_OFN1_TL02_PHS0_sel_0, Z => TL02_kb_y_6);
  g672 : AO22D0BWP7T port map(A1 => diry1new2(4), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => diry2new2(4), Z => TL02_kb_y_4);
  g673 : AO22D0BWP7T port map(A1 => diry1new2(1), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => diry2new2(1), Z => TL02_kb_y_1);
  g676 : AO32D0BWP7T port map(A1 => n_479, A2 => FE_PHN174_vcountintern_8, A3 => FE_DBTN14_reset, B1 => vcountintern(9), B2 => FE_DBTN14_reset, Z => n_480);
  g677 : ND2D1BWP7T port map(A1 => n_478, A2 => n_508, ZN => n_479);
  g678 : AOI31D0BWP7T port map(A1 => vcountintern(2), A2 => vcountintern(1), A3 => vcountintern(0), B => vcountintern(3), ZN => n_478);
  buf4_stored_reg_7 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_17, D => diry1new1(7), Q => diry1new2(7));
  buf3_stored_reg_4 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_17, D => dirx1new1(4), Q => dirx1new2(4));
  buf5_stored_reg_3 : DFKCNQD1BWP7T port map(CN => TL01_n_63, CP => CTS_17, D => dirx2new1(3), Q => dirx2new2(3));
  buf3_stored_reg_3 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_17, D => dirx1new1(3), Q => dirx1new2(3));
  buf5_stored_reg_2 : DFKCNQD1BWP7T port map(CN => TL01_n_63, CP => CTS_17, D => dirx2new1(2), Q => dirx2new2(2));
  buf3_stored_reg_2 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_17, D => dirx1new1(2), Q => dirx1new2(2));
  buf5_stored_reg_1 : DFKCNQD1BWP7T port map(CN => TL01_n_63, CP => CTS_17, D => dirx2new1(1), Q => dirx2new2(1));
  buf6_stored_reg_7 : DFKCNQD1BWP7T port map(CN => diry2new1(7), CP => CTS_17, D => TL01_n_63, Q => diry2new2(7));
  buf5_stored_reg_4 : DFKCNQD1BWP7T port map(CN => TL01_n_63, CP => CTS_17, D => dirx2new1(4), Q => dirx2new2(4));
  buf4_stored_reg_6 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_17, D => diry1new1(6), Q => diry1new2(6));
  buf5_stored_reg_7 : DFKCNQD1BWP7T port map(CN => TL01_n_63, CP => CTS_17, D => dirx2new1(7), Q => dirx2new2(7));
  buf6_stored_reg_5 : DFKCNQD1BWP7T port map(CN => TL01_n_63, CP => CTS_17, D => diry2new1(5), Q => diry2new2(5));
  buf3_stored_reg_7 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_17, D => dirx1new1(7), Q => dirx1new2(7));
  buf3_stored_reg_5 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_17, D => dirx1new1(5), Q => dirx1new2(5));
  buf5_stored_reg_6 : DFKCNQD1BWP7T port map(CN => TL01_n_63, CP => CTS_17, D => dirx2new1(6), Q => dirx2new2(6));
  buf6_stored_reg_6 : DFKCNQD1BWP7T port map(CN => TL01_n_63, CP => CTS_17, D => diry2new1(6), Q => diry2new2(6));
  buf5_stored_reg_5 : DFKCNQD1BWP7T port map(CN => TL01_n_63, CP => CTS_17, D => dirx2new1(5), Q => dirx2new2(5));
  buf3_stored_reg_6 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_17, D => dirx1new1(6), Q => dirx1new2(6));
  TL00_DM10_mem_reg_0_0 : DFQD1BWP7T port map(CP => CTS_17, D => n_110, Q => char1perc(0));
  TL00_DM10_mem_reg_0_1 : DFQD1BWP7T port map(CP => CTS_17, D => n_102, Q => char1perc(1));
  TL00_DM10_mem_reg_0_2 : DFQD1BWP7T port map(CP => CTS_17, D => n_100, Q => char1perc(2));
  TL00_DM10_mem_reg_0_3 : DFQD1BWP7T port map(CP => CTS_17, D => n_97, Q => char1perc(3));
  TL00_DM10_mem_reg_0_4 : DFQD1BWP7T port map(CP => CTS_17, D => n_114, Q => char1perc(4));
  TL00_DM10_mem_reg_0_5 : DFQD1BWP7T port map(CP => CTS_17, D => n_96, Q => char1perc(5));
  TL00_DM10_mem_reg_0_6 : DFQD1BWP7T port map(CP => CTS_17, D => n_95, Q => char1perc(6));
  TL00_DM10_mem_reg_0_7 : DFQD1BWP7T port map(CP => CTS_17, D => n_94, Q => char1perc(7));
  TL00_DM11_mem_reg_0_0 : DFQD1BWP7T port map(CP => CTS_17, D => n_93, Q => char2perc(0));
  TL00_DM11_mem_reg_0_1 : DFQD1BWP7T port map(CP => CTS_17, D => n_106, Q => char2perc(1));
  TL00_DM11_mem_reg_0_2 : DFQD1BWP7T port map(CP => CTS_17, D => n_92, Q => char2perc(2));
  TL00_DM11_mem_reg_0_3 : DFQD1BWP7T port map(CP => CTS_17, D => n_103, Q => char2perc(3));
  TL00_DM11_mem_reg_0_4 : DFQD1BWP7T port map(CP => CTS_17, D => n_104, Q => char2perc(4));
  TL00_DM11_mem_reg_0_5 : DFQD1BWP7T port map(CP => CTS_17, D => n_91, Q => char2perc(5));
  TL00_DM11_mem_reg_0_6 : DFQD1BWP7T port map(CP => CTS_17, D => n_90, Q => char2perc(6));
  TL00_DM11_mem_reg_0_7 : DFQD1BWP7T port map(CP => CTS_17, D => n_89, Q => char2perc(7));
  TL00_DM20_mem_reg_0_0 : DFQD1BWP7T port map(CP => CTS_16, D => FE_PHN127_n_88, Q => char1posx(0));
  TL00_DM20_mem_reg_0_1 : DFQD1BWP7T port map(CP => CTS_15, D => FE_PHN132_n_75, Q => char1posx(1));
  TL00_DM20_mem_reg_0_2 : DFQD1BWP7T port map(CP => CTS_15, D => FE_PHN134_n_72, Q => char1posx(2));
  TL00_DM20_mem_reg_0_3 : DFQD1BWP7T port map(CP => CTS_16, D => FE_PHN130_n_98, Q => char1posx(3));
  TL00_DM20_mem_reg_0_4 : DFQD1BWP7T port map(CP => CTS_15, D => FE_PHN128_n_113, Q => char1posx(4));
  TL00_DM20_mem_reg_0_5 : DFQD1BWP7T port map(CP => CTS_15, D => n_101, Q => char1posx(5));
  TL00_DM20_mem_reg_0_6 : DFQD1BWP7T port map(CP => CTS_15, D => FE_PHN133_n_70, Q => char1posx(6));
  TL00_DM20_mem_reg_0_7 : DFQD1BWP7T port map(CP => CTS_15, D => FE_PHN141_n_109, Q => char1posx(7));
  TL00_DM20_mem_reg_0_8 : DFQD1BWP7T port map(CP => CTS_15, D => n_112, Q => FE_PHN124_char1posx_8);
  TL00_DM21_mem_reg_0_0 : DFQD1BWP7T port map(CP => CTS_17, D => FE_PHN137_n_111, Q => char1posy(0));
  TL00_DM21_mem_reg_0_1 : DFQD1BWP7T port map(CP => CTS_17, D => FE_PHN142_n_108, Q => char1posy(1));
  TL00_DM21_mem_reg_0_2 : DFQD1BWP7T port map(CP => CTS_16, D => n_71, Q => char1posy(2));
  TL00_DM21_mem_reg_0_3 : DFQD1BWP7T port map(CP => CTS_17, D => n_107, Q => char1posy(3));
  TL00_DM21_mem_reg_0_4 : DFQD1BWP7T port map(CP => CTS_17, D => FE_PHN131_n_105, Q => char1posy(4));
  TL00_DM21_mem_reg_0_5 : DFQD1BWP7T port map(CP => CTS_15, D => FE_PHN139_n_74, Q => char1posy(5));
  TL00_DM21_mem_reg_0_6 : DFQD1BWP7T port map(CP => CTS_16, D => n_73, Q => char1posy(6));
  TL00_DM21_mem_reg_0_7 : DFQD1BWP7T port map(CP => CTS_17, D => FE_PHN135_n_99, Q => char1posy(7));
  TL00_DM22_mem_reg_0_0 : DFQD1BWP7T port map(CP => CTS_15, D => n_350, Q => char2posx(0));
  TL00_DM22_mem_reg_0_1 : DFQD1BWP7T port map(CP => CTS_15, D => n_356, Q => char2posx(1));
  TL00_DM22_mem_reg_0_2 : DFQD1BWP7T port map(CP => CTS_15, D => n_361, Q => char2posx(2));
  TL00_DM22_mem_reg_0_3 : DFQD1BWP7T port map(CP => CTS_15, D => n_367, Q => char2posx(3));
  TL00_DM22_mem_reg_0_4 : DFQD1BWP7T port map(CP => CTS_15, D => n_375, Q => char2posx(4));
  TL00_DM22_mem_reg_0_5 : DFQD1BWP7T port map(CP => CTS_15, D => n_385, Q => char2posx(5));
  TL00_DM22_mem_reg_0_6 : DFQD1BWP7T port map(CP => CTS_15, D => n_399, Q => char2posx(6));
  TL00_DM22_mem_reg_0_7 : DFQD1BWP7T port map(CP => CTS_15, D => n_411, Q => char2posx(7));
  TL00_DM22_mem_reg_0_8 : DFQD1BWP7T port map(CP => CTS_15, D => n_414, Q => char2posx(8));
  TL00_DM23_mem_reg_0_0 : DFQD1BWP7T port map(CP => CTS_17, D => n_435, Q => char2posy(0));
  TL00_DM23_mem_reg_0_1 : DFQD1BWP7T port map(CP => CTS_17, D => n_462, Q => char2posy(1));
  TL00_DM23_mem_reg_0_2 : DFQD1BWP7T port map(CP => CTS_16, D => n_474, Q => char2posy(2));
  TL00_DM23_mem_reg_0_3 : DFQD1BWP7T port map(CP => CTS_17, D => n_469, Q => char2posy(3));
  TL00_DM23_mem_reg_0_4 : DFQD1BWP7T port map(CP => CTS_17, D => n_468, Q => char2posy(4));
  TL00_DM23_mem_reg_0_5 : DFQD1BWP7T port map(CP => CTS_17, D => n_472, Q => char2posy(5));
  TL00_DM23_mem_reg_0_6 : DFQD1BWP7T port map(CP => CTS_17, D => n_456, Q => char2posy(6));
  TL00_DM23_mem_reg_0_7 : DFQD1BWP7T port map(CP => CTS_17, D => n_265, Q => char2posy(7));
  TL00_DM30_mem_reg_0_0 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_15, D => FE_PHN32_char1velxin_0, E => FE_OFN4_TL00_writeint, Q => char1velx(0));
  TL00_DM30_mem_reg_0_1 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_15, D => char1velxin(1), E => FE_OFN4_TL00_writeint, Q => char1velx(1));
  TL00_DM30_mem_reg_0_2 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_15, D => FE_PHN25_char1velxin_2, E => FE_OFN4_TL00_writeint, Q => char1velx(2));
  TL00_DM30_mem_reg_0_3 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_15, D => char1velxin(3), E => FE_OFN4_TL00_writeint, Q => char1velx(3));
  TL00_DM30_mem_reg_0_4 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_15, D => FE_PHN22_char1velxin_4, E => FE_OFN4_TL00_writeint, Q => char1velx(4));
  TL00_DM30_mem_reg_0_5 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_15, D => FE_PHN27_char1velxin_5, E => FE_OFN4_TL00_writeint, Q => char1velx(5));
  TL00_DM30_mem_reg_0_6 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_17, D => char1velxin(6), E => FE_OFN4_TL00_writeint, Q => char1velx(6));
  TL00_DM30_mem_reg_0_7 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_15, D => char1velxin(7), E => FE_OFN4_TL00_writeint, Q => char1velx(7));
  TL00_DM30_mem_reg_0_8 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_15, D => FE_PHN61_char1velxin_8, E => FE_OFN4_TL00_writeint, Q => char1velx(8));
  TL00_DM30_mem_reg_0_9 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_15, D => FE_PHN21_char1velxin_9, E => FE_OFN4_TL00_writeint, Q => char1velx(9));
  TL00_DM31_mem_reg_0_0 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_17, D => char1velyin(0), E => FE_OFN4_TL00_writeint, Q => char1vely(0));
  TL00_DM31_mem_reg_0_1 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_17, D => char1velyin(1), E => FE_OFN4_TL00_writeint, Q => char1vely(1));
  TL00_DM31_mem_reg_0_2 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_15, D => FE_PHN30_char1velyin_2, E => FE_OFN4_TL00_writeint, Q => char1vely(2));
  TL00_DM31_mem_reg_0_3 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_15, D => FE_PHN24_char1velyin_3, E => FE_OFN4_TL00_writeint, Q => char1vely(3));
  TL00_DM31_mem_reg_0_4 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_17, D => FE_PHN31_char1velyin_4, E => FE_OFN4_TL00_writeint, Q => char1vely(4));
  TL00_DM31_mem_reg_0_5 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_15, D => char1velyin(5), E => FE_OFN4_TL00_writeint, Q => char1vely(5));
  TL00_DM31_mem_reg_0_6 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_15, D => FE_PHN39_char1velyin_6, E => FE_OFN4_TL00_writeint, Q => char1vely(6));
  TL00_DM31_mem_reg_0_7 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_15, D => char1velyin(7), E => FE_OFN4_TL00_writeint, Q => char1vely(7));
  TL00_DM31_mem_reg_0_8 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_17, D => char1velyin(8), E => FE_OFN4_TL00_writeint, Q => char1vely(8));
  TL00_DM31_mem_reg_0_9 : EDFKCNQD1BWP7T port map(CN => n_16, CP => CTS_17, D => char1velyin(9), E => FE_OFN4_TL00_writeint, Q => char1vely(9));
  TL00_DM32_mem_reg_0_0 : DFKCNQD1BWP7T port map(CN => n_13, CP => CTS_15, D => n_326, Q => char2velx(0));
  TL00_DM32_mem_reg_0_1 : DFKCNQD1BWP7T port map(CN => n_13, CP => CTS_15, D => n_348, Q => char2velx(1));
  TL00_DM32_mem_reg_0_2 : DFKCNQD1BWP7T port map(CN => n_13, CP => CTS_15, D => n_341, Q => char2velx(2));
  TL00_DM32_mem_reg_0_3 : DFKCNQD1BWP7T port map(CN => n_13, CP => CTS_15, D => n_336, Q => char2velx(3));
  TL00_DM32_mem_reg_0_4 : DFKCNQD1BWP7T port map(CN => n_13, CP => CTS_15, D => n_346, Q => char2velx(4));
  TL00_DM32_mem_reg_0_5 : DFKCNQD1BWP7T port map(CN => n_13, CP => CTS_15, D => n_339, Q => char2velx(5));
  TL00_DM32_mem_reg_0_6 : EDFKCNQD1BWP7T port map(CN => n_13, CP => CTS_15, D => n_320, E => FE_OFN4_TL00_writeint, Q => char2velx(6));
  TL00_DM32_mem_reg_0_7 : DFKCNQD1BWP7T port map(CN => n_13, CP => CTS_15, D => n_334, Q => char2velx(7));
  TL00_DM32_mem_reg_0_8 : EDFKCNQD1BWP7T port map(CN => n_13, CP => CTS_15, D => n_324, E => FE_OFN4_TL00_writeint, Q => char2velx(8));
  TL00_DM32_mem_reg_0_9 : DFKCNQD1BWP7T port map(CN => n_13, CP => CTS_15, D => n_333, Q => char2velx(9));
  TL00_DM33_mem_reg_0_0 : EDFKCNQD1BWP7T port map(CN => n_13, CP => CTS_15, D => n_451, E => FE_OFN4_TL00_writeint, Q => char2vely(0));
  TL00_DM33_mem_reg_0_1 : EDFKCNQD1BWP7T port map(CN => n_13, CP => CTS_17, D => n_444, E => FE_OFN4_TL00_writeint, Q => char2vely(1));
  TL00_DM33_mem_reg_0_2 : EDFKCNQD1BWP7T port map(CN => n_13, CP => CTS_17, D => n_443, E => FE_OFN4_TL00_writeint, Q => char2vely(2));
  TL00_DM33_mem_reg_0_3 : DFKCNQD1BWP7T port map(CN => n_13, CP => CTS_15, D => n_453, Q => FE_PHN175_char2vely_3);
  TL00_DM33_mem_reg_0_4 : EDFKCNQD1BWP7T port map(CN => n_13, CP => CTS_17, D => n_442, E => FE_OFN4_TL00_writeint, Q => char2vely(4));
  TL00_DM33_mem_reg_0_5 : EDFKCNQD1BWP7T port map(CN => n_13, CP => CTS_15, D => n_440, E => FE_OFN4_TL00_writeint, Q => char2vely(5));
  TL00_DM33_mem_reg_0_6 : EDFKCNQD1BWP7T port map(CN => n_13, CP => CTS_15, D => n_438, E => FE_OFN4_TL00_writeint, Q => char2vely(6));
  TL00_DM33_mem_reg_0_7 : EDFKCNQD1BWP7T port map(CN => n_13, CP => CTS_17, D => n_437, E => FE_OFN4_TL00_writeint, Q => char2vely(7));
  TL00_DM33_mem_reg_0_8 : EDFKCNQD1BWP7T port map(CN => n_13, CP => CTS_17, D => n_441, E => FE_OFN4_TL00_writeint, Q => char2vely(8));
  TL00_DM33_mem_reg_0_9 : EDFKCNQD1BWP7T port map(CN => n_13, CP => CTS_17, D => n_439, E => FE_OFN4_TL00_writeint, Q => char2vely(9));
  TL00_WL00_state_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => n_56, Q => TL00_WL00_state_1);
  TL02_PHS0_px1m_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => n_351, Q => FE_PHN49_char1posxin_0);
  TL02_PHS0_px1m_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_15, D => n_355, Q => char1posxin(1));
  TL02_PHS0_px1m_reg_2 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_15, D => n_360, Q => FE_PHN56_char1posxin_2);
  TL02_PHS0_px1m_reg_3 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => n_366, Q => char1posxin(3));
  TL02_PHS0_px1m_reg_4 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_15, D => n_371, Q => char1posxin(4));
  TL02_PHS0_px1m_reg_5 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_15, D => n_380, Q => char1posxin(5));
  TL02_PHS0_px1m_reg_6 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_15, D => n_393, Q => char1posxin(6));
  TL02_PHS0_px1m_reg_7 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_15, D => n_404, Q => FE_PHN57_char1posxin_7);
  TL02_PHS0_px1m_reg_8 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_15, D => n_415, Q => char1posxin(8));
  TL02_PHS0_py1m_reg_0 : DFQD1BWP7T port map(CP => CTS_15, D => n_454, Q => FE_PHN41_char1posyin_0);
  TL02_PHS0_py1m_reg_1 : DFQD1BWP7T port map(CP => CTS_15, D => n_473, Q => FE_PHN63_char1posyin_1);
  TL02_PHS0_py1m_reg_2 : DFQD1BWP7T port map(CP => CTS_15, D => n_457, Q => FE_PHN47_char1posyin_2);
  TL02_PHS0_py1m_reg_3 : DFQD1BWP7T port map(CP => CTS_17, D => n_471, Q => FE_PHN44_char1posyin_3);
  TL02_PHS0_py1m_reg_4 : DFQD1BWP7T port map(CP => CTS_17, D => n_470, Q => FE_PHN42_char1posyin_4);
  TL02_PHS0_py1m_reg_5 : DFQD1BWP7T port map(CP => CTS_15, D => n_455, Q => FE_PHN43_char1posyin_5);
  TL02_PHS0_py1m_reg_6 : DFQD1BWP7T port map(CP => CTS_17, D => n_434, Q => FE_PHN45_char1posyin_6);
  TL02_PHS0_py1m_reg_7 : DFQD1BWP7T port map(CP => CTS_17, D => n_266, Q => char1posyin(7));
  TL02_PHS0_vx1m_reg_0 : DFQD1BWP7T port map(CP => CTS_15, D => n_327, Q => char1velxin(0));
  TL02_PHS0_vx1m_reg_1 : DFQD1BWP7T port map(CP => CTS_15, D => n_349, Q => FE_PHN29_char1velxin_1);
  TL02_PHS0_vx1m_reg_2 : DFQD1BWP7T port map(CP => CTS_15, D => n_345, Q => char1velxin(2));
  TL02_PHS0_vx1m_reg_3 : DFQD1BWP7T port map(CP => CTS_15, D => n_332, Q => FE_PHN26_char1velxin_3);
  TL02_PHS0_vx1m_reg_4 : DFQD1BWP7T port map(CP => CTS_15, D => n_342, Q => char1velxin(4));
  TL02_PHS0_vx1m_reg_5 : DFQD1BWP7T port map(CP => CTS_15, D => n_335, Q => char1velxin(5));
  TL02_PHS0_vx1m_reg_6 : DFQD1BWP7T port map(CP => CTS_15, D => n_344, Q => FE_PHN36_char1velxin_6);
  TL02_PHS0_vx1m_reg_7 : DFQD1BWP7T port map(CP => CTS_15, D => n_338, Q => FE_PHN23_char1velxin_7);
  TL02_PHS0_vx1m_reg_8 : DFQD1BWP7T port map(CP => CTS_17, D => n_343, Q => char1velxin(8));
  TL02_PHS0_vx1m_reg_9 : DFQD1BWP7T port map(CP => CTS_15, D => n_337, Q => char1velxin(9));
  TL02_PHS0_vy1m_reg_0 : DFQD1BWP7T port map(CP => CTS_15, D => n_461, Q => FE_PHN33_char1velyin_0);
  TL02_PHS0_vy1m_reg_1 : DFQD1BWP7T port map(CP => CTS_17, D => n_465, Q => FE_PHN35_char1velyin_1);
  TL02_PHS0_vy1m_reg_2 : DFQD1BWP7T port map(CP => CTS_17, D => n_466, Q => char1velyin(2));
  TL02_PHS0_vy1m_reg_3 : DFQD1BWP7T port map(CP => CTS_15, D => n_452, Q => char1velyin(3));
  TL02_PHS0_vy1m_reg_4 : DFQD1BWP7T port map(CP => CTS_15, D => n_464, Q => char1velyin(4));
  TL02_PHS0_vy1m_reg_5 : DFQD1BWP7T port map(CP => CTS_15, D => n_463, Q => FE_PHN28_char1velyin_5);
  TL02_PHS0_vy1m_reg_6 : DFQD1BWP7T port map(CP => CTS_15, D => n_467, Q => char1velyin(6));
  TL02_PHS0_vy1m_reg_7 : DFQD1BWP7T port map(CP => CTS_15, D => n_460, Q => FE_PHN37_char1velyin_7);
  TL02_PHS0_vy1m_reg_8 : DFQD1BWP7T port map(CP => CTS_17, D => n_458, Q => FE_PHN38_char1velyin_8);
  TL02_PHS0_vy1m_reg_9 : DFQD1BWP7T port map(CP => CTS_17, D => n_459, Q => FE_PHN40_char1velyin_9);
  buf3_stored_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_17, D => dirx1new1(0), Q => dirx1new2(0));
  buf3_stored_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_17, D => dirx1new1(1), Q => dirx1new2(1));
  buf4_stored_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_17, D => diry1new1(0), Q => diry1new2(0));
  buf4_stored_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_17, D => diry1new1(1), Q => diry1new2(1));
  buf4_stored_reg_2 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_17, D => diry1new1(2), Q => diry1new2(2));
  buf4_stored_reg_3 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_17, D => diry1new1(3), Q => diry1new2(3));
  buf4_stored_reg_4 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_17, D => diry1new1(4), Q => diry1new2(4));
  buf4_stored_reg_5 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_17, D => diry1new1(5), Q => diry1new2(5));
  buf5_stored_reg_0 : DFKCNQD1BWP7T port map(CN => TL01_n_63, CP => CTS_17, D => dirx2new1(0), Q => dirx2new2(0));
  buf6_stored_reg_0 : DFKCNQD1BWP7T port map(CN => TL01_n_63, CP => CTS_17, D => diry2new1(0), Q => diry2new2(0));
  buf6_stored_reg_1 : DFKCNQD1BWP7T port map(CN => TL01_n_63, CP => CTS_17, D => diry2new1(1), Q => diry2new2(1));
  buf6_stored_reg_2 : DFKCNQD1BWP7T port map(CN => TL01_n_63, CP => CTS_17, D => diry2new1(2), Q => diry2new2(2));
  buf6_stored_reg_3 : DFKCNQD1BWP7T port map(CN => TL01_n_63, CP => CTS_17, D => diry2new1(3), Q => diry2new2(3));
  buf6_stored_reg_4 : DFKCNQD1BWP7T port map(CN => TL01_n_63, CP => CTS_17, D => diry2new1(4), Q => diry2new2(4));
  g7085 : AO221D0BWP7T port map(A1 => n_445, A2 => FE_OFN4_TL00_writeint, B1 => n_1, B2 => FE_PHN101_char2posy_2, C => n_12, Z => n_474);
  g7095 : MOAI22D0BWP7T port map(A1 => n_446, A2 => n_136, B1 => n_135, B2 => FE_PHN177_char1posyin_1, ZN => n_473);
  g7096 : AO211D0BWP7T port map(A1 => n_1, A2 => FE_PHN72_char2posy_5, B => n_436, C => n_12, Z => n_472);
  g7097 : AO22D0BWP7T port map(A1 => n_449, A2 => n_137, B1 => char1posyin(3), B2 => n_135, Z => n_471);
  g7098 : AO22D0BWP7T port map(A1 => n_447, A2 => n_137, B1 => char1posyin(4), B2 => n_135, Z => n_470);
  g7099 : MOAI22D0BWP7T port map(A1 => n_450, A2 => n_59, B1 => n_61, B2 => FE_PHN83_char2posy_3, ZN => n_469);
  g7100 : MOAI22D0BWP7T port map(A1 => n_448, A2 => n_59, B1 => n_61, B2 => FE_PHN79_char2posy_4, ZN => n_468);
  g7105 : AO22D0BWP7T port map(A1 => n_438, A2 => n_137, B1 => FE_PHN39_char1velyin_6, B2 => n_135, Z => n_467);
  g7106 : AO22D0BWP7T port map(A1 => n_443, A2 => n_137, B1 => FE_PHN30_char1velyin_2, B2 => n_135, Z => n_466);
  g7107 : AO22D0BWP7T port map(A1 => n_444, A2 => n_137, B1 => char1velyin(1), B2 => n_135, Z => n_465);
  g7108 : AO22D0BWP7T port map(A1 => n_442, A2 => n_137, B1 => FE_PHN31_char1velyin_4, B2 => n_135, Z => n_464);
  g7109 : AO22D0BWP7T port map(A1 => n_440, A2 => n_137, B1 => char1velyin(5), B2 => n_135, Z => n_463);
  g7110 : MOAI22D0BWP7T port map(A1 => n_446, A2 => n_59, B1 => n_61, B2 => FE_PHN81_char2posy_1, ZN => n_462);
  g7111 : AO22D0BWP7T port map(A1 => n_451, A2 => n_137, B1 => char1velyin(0), B2 => n_135, Z => n_461);
  g7112 : AO22D0BWP7T port map(A1 => n_437, A2 => n_137, B1 => char1velyin(7), B2 => n_135, Z => n_460);
  g7113 : AO22D0BWP7T port map(A1 => n_439, A2 => n_137, B1 => char1velyin(9), B2 => n_135, Z => n_459);
  g7114 : AO22D0BWP7T port map(A1 => n_441, A2 => n_137, B1 => char1velyin(8), B2 => n_135, Z => n_458);
  g7115 : AO22D0BWP7T port map(A1 => n_445, A2 => n_137, B1 => char1posyin(2), B2 => n_135, Z => n_457);
  g7116 : AO221D0BWP7T port map(A1 => n_431, A2 => FE_OFN4_TL00_writeint, B1 => n_1, B2 => FE_PHN93_char2posy_6, C => n_12, Z => n_456);
  g7119 : MOAI22D0BWP7T port map(A1 => n_0, A2 => n_230, B1 => n_135, B2 => char1posyin(5), ZN => n_455);
  g7120 : MOAI22D0BWP7T port map(A1 => n_0, A2 => n_139, B1 => n_135, B2 => char1posyin(0), ZN => n_454);
  g7121 : OAI31D0BWP7T port map(A1 => n_1, A2 => n_164, A3 => n_432, B => n_11, ZN => n_453);
  g7122 : MOAI22D0BWP7T port map(A1 => n_0, A2 => n_164, B1 => n_135, B2 => FE_PHN24_char1velyin_3, ZN => n_452);
  g7123 : INVD0BWP7T port map(I => n_449, ZN => n_450);
  g7124 : INVD0BWP7T port map(I => n_447, ZN => n_448);
  g7125 : OAI21D0BWP7T port map(A1 => n_432, A2 => n_115, B => n_433, ZN => n_451);
  g7126 : OAI21D0BWP7T port map(A1 => n_432, A2 => n_198, B => n_430, ZN => n_449);
  g7127 : OAI21D0BWP7T port map(A1 => n_432, A2 => n_214, B => n_428, ZN => n_447);
  g7128 : OA21D0BWP7T port map(A1 => n_432, A2 => n_162, B => n_430, Z => n_446);
  g7129 : OAI21D0BWP7T port map(A1 => n_432, A2 => n_183, B => n_429, ZN => n_445);
  g7130 : OAI21D0BWP7T port map(A1 => n_432, A2 => n_138, B => n_433, ZN => n_444);
  g7131 : OAI21D0BWP7T port map(A1 => n_432, A2 => n_147, B => n_433, ZN => n_443);
  g7132 : OAI21D0BWP7T port map(A1 => n_432, A2 => n_169, B => n_433, ZN => n_442);
  g7133 : NR3D0BWP7T port map(A1 => n_432, A2 => n_230, A3 => n_1, ZN => n_436);
  g7134 : OAI31D0BWP7T port map(A1 => n_59, A2 => n_139, A3 => n_432, B => n_78, ZN => n_435);
  g7135 : AO22D0BWP7T port map(A1 => n_431, A2 => n_137, B1 => char1posyin(6), B2 => n_135, Z => n_434);
  g7136 : OAI21D0BWP7T port map(A1 => n_432, A2 => n_237, B => n_433, ZN => n_441);
  g7137 : OAI21D0BWP7T port map(A1 => n_432, A2 => n_174, B => n_433, ZN => n_440);
  g7138 : OAI21D0BWP7T port map(A1 => n_432, A2 => n_253, B => n_433, ZN => n_439);
  g7139 : OAI21D0BWP7T port map(A1 => n_432, A2 => n_205, B => n_433, ZN => n_438);
  g7140 : OAI21D0BWP7T port map(A1 => n_432, A2 => n_216, B => n_433, ZN => n_437);
  g7142 : OAI221D1BWP7T port map(A1 => inputsp1(2), A2 => FE_OFN1_TL02_PHS0_sel_0, B1 => FE_OFN0_n_6, B2 => inputsp2(2), C => n_432, ZN => n_433);
  g7144 : ND2D1BWP7T port map(A1 => n_430, A2 => n_428, ZN => n_432);
  g7145 : ND2D1BWP7T port map(A1 => n_430, A2 => n_236, ZN => n_431);
  g7146 : OA211D0BWP7T port map(A1 => n_236, A2 => n_254, B => n_429, C => n_252, Z => n_430);
  g7147 : OR4D1BWP7T port map(A1 => n_236, A2 => n_263, A3 => n_262, A4 => n_427, Z => n_429);
  g7148 : ND4D0BWP7T port map(A1 => n_426, A2 => n_252, A3 => n_243, A4 => n_236, ZN => n_428);
  g7149 : OAI211D1BWP7T port map(A1 => n_251, A2 => n_255, B => n_425, C => n_264, ZN => n_427);
  g7150 : NR2XD0BWP7T port map(A1 => n_424, A2 => n_263, ZN => n_426);
  g7151 : OAI31D0BWP7T port map(A1 => n_406, A2 => n_390, A3 => n_407, B => n_423, ZN => n_425);
  g7152 : OAI222D0BWP7T port map(A1 => n_248, A2 => n_251, B1 => n_162, B2 => n_264, C1 => n_418, C2 => n_422, ZN => n_424);
  g7153 : AOI33D1BWP7T port map(A1 => n_417, A2 => n_364, A3 => n_358, B1 => n_421, B2 => n_401, B3 => n_353, ZN => n_423);
  g7154 : OAI211D1BWP7T port map(A1 => n_416, A2 => n_419, B => n_420, C => n_413, ZN => n_422);
  g7156 : NR3D0BWP7T port map(A1 => n_416, A2 => n_387, A3 => n_365, ZN => n_421);
  g7158 : OAI21D0BWP7T port map(A1 => n_410, A2 => n_409, B => n_416, ZN => n_420);
  g7159 : AOI221D0BWP7T port map(A1 => n_410, A2 => n_378, B1 => n_397, B2 => n_379, C => n_408, ZN => n_419);
  g7160 : AOI211XD0BWP7T port map(A1 => n_382, A2 => n_389, B => n_412, C => n_376, ZN => n_418);
  g7161 : AOI211XD0BWP7T port map(A1 => n_353, A2 => n_328, B => n_412, C => n_391, ZN => n_417);
  g7164 : MOAI22D0BWP7T port map(A1 => n_405, A2 => n_127, B1 => n_127, B2 => FE_PHN52_char1posxin_8, ZN => n_415);
  g7165 : MOAI22D0BWP7T port map(A1 => n_405, A2 => n_59, B1 => n_61, B2 => FE_PHN123_char2posx_8, ZN => n_414);
  g7166 : OR3D1BWP7T port map(A1 => n_389, A2 => n_406, A3 => n_396, Z => n_413);
  g7167 : MOAI22D0BWP7T port map(A1 => n_402, A2 => n_406, B1 => n_402, B2 => n_406, ZN => n_416);
  g7168 : ND2D1BWP7T port map(A1 => n_407, A2 => n_405, ZN => n_412);
  g7169 : AO221D0BWP7T port map(A1 => n_401, A2 => FE_OFN4_TL00_writeint, B1 => n_1, B2 => char2posx(7), C => n_12, Z => n_411);
  g7170 : AOI21D0BWP7T port map(A1 => n_387, A2 => n_358, B => n_403, ZN => n_409);
  g7171 : NR4D0BWP7T port map(A1 => n_397, A2 => n_400, A3 => n_379, A4 => n_364, ZN => n_408);
  g7172 : NR2D1BWP7T port map(A1 => n_403, A2 => n_364, ZN => n_410);
  g7173 : INVD0BWP7T port map(I => n_406, ZN => n_405);
  g7174 : MOAI22D0BWP7T port map(A1 => n_400, A2 => n_127, B1 => n_127, B2 => char1posxin(7), ZN => n_404);
  g7175 : MAOI22D0BWP7T port map(A1 => n_400, A2 => n_398, B1 => n_400, B2 => n_398, ZN => n_407);
  g7176 : MOAI22D0BWP7T port map(A1 => n_395, A2 => n_340, B1 => n_395, B2 => n_340, ZN => n_406);
  g7177 : OR2D1BWP7T port map(A1 => n_397, A2 => n_401, Z => n_403);
  g7178 : ND2D1BWP7T port map(A1 => n_400, A2 => n_392, ZN => n_402);
  g7179 : INVD1BWP7T port map(I => n_400, ZN => n_401);
  g7182 : MAOI22D0BWP7T port map(A1 => n_504, A2 => n_30, B1 => n_504, B2 => n_30, ZN => n_400);
  g7183 : AO221D0BWP7T port map(A1 => n_381, A2 => FE_OFN4_TL00_writeint, B1 => n_1, B2 => FE_PHN119_char2posx_6, C => n_12, Z => n_399);
  g7184 : OAI211D1BWP7T port map(A1 => n_354, A2 => n_364, B => n_386, C => n_365, ZN => n_396);
  g7185 : NR3D0BWP7T port map(A1 => n_377, A2 => n_389, A3 => n_364, ZN => n_398);
  g7186 : AO21D0BWP7T port map(A1 => n_384, A2 => n_381, B => n_392, Z => n_397);
  g7187 : MOAI22D0BWP7T port map(A1 => n_389, A2 => n_127, B1 => n_127, B2 => FE_PHN162_char1posxin_6, ZN => n_393);
  g7188 : MAOI222D1BWP7T port map(A => n_383, B => n_318, C => n_30, ZN => n_395);
  g7192 : INVD0BWP7T port map(I => n_390, ZN => n_391);
  g7193 : NR2XD0BWP7T port map(A1 => n_384, A2 => n_381, ZN => n_392);
  g7194 : NR3D0BWP7T port map(A1 => n_382, A2 => n_373, A3 => n_389, ZN => n_390);
  g7195 : INVD1BWP7T port map(I => n_381, ZN => n_389);
  g7197 : INVD0BWP7T port map(I => n_386, ZN => n_387);
  g7198 : ND2D1BWP7T port map(A1 => n_382, A2 => n_373, ZN => n_386);
  g7199 : AO221D0BWP7T port map(A1 => n_378, A2 => FE_OFN4_TL00_writeint, B1 => n_1, B2 => char2posx(5), C => n_12, Z => n_385);
  g7200 : ND3D0BWP7T port map(A1 => n_377, A2 => n_369, A3 => n_364, ZN => n_384);
  g7201 : AOI21D0BWP7T port map(A1 => n_374, A2 => n_330, B => n_331, ZN => n_383);
  g7202 : MOAI22D0BWP7T port map(A1 => n_377, A2 => n_127, B1 => n_127, B2 => FE_PHN167_char1posxin_5, ZN => n_380);
  g7203 : MAOI22D0BWP7T port map(A1 => n_377, A2 => n_370, B1 => n_377, B2 => n_370, ZN => n_382);
  g7204 : MOAI22D0BWP7T port map(A1 => n_374, A2 => n_347, B1 => n_374, B2 => n_347, ZN => n_381);
  g7205 : OR2D1BWP7T port map(A1 => n_373, A2 => n_378, Z => n_379);
  g7206 : INVD0BWP7T port map(I => n_377, ZN => n_378);
  g7209 : INR3D0BWP7T port map(A1 => n_373, B1 => n_354, B2 => n_365, ZN => n_376);
  g7210 : MAOI22D0BWP7T port map(A1 => n_372, A2 => n_323, B1 => n_372, B2 => n_323, ZN => n_377);
  g7211 : OAI211D1BWP7T port map(A1 => n_1, A2 => n_369, B => n_13, C => n_14, ZN => n_375);
  g7212 : MAOI222D1BWP7T port map(A => n_368, B => n_323, C => n_62, ZN => n_374);
  g7213 : MAOI22D0BWP7T port map(A1 => n_369, A2 => n_363, B1 => n_369, B2 => n_363, ZN => n_373);
  g7214 : MOAI22D0BWP7T port map(A1 => n_369, A2 => n_127, B1 => n_127, B2 => FE_PHN50_char1posxin_4, ZN => n_371);
  g7215 : CKXOR2D1BWP7T port map(A1 => n_368, A2 => n_62, Z => n_372);
  g7216 : NR2D1BWP7T port map(A1 => n_369, A2 => n_364, ZN => n_370);
  g7217 : FA1D0BWP7T port map(A => n_317, B => n_51, CI => n_362, CO => n_368, S => n_369);
  g7220 : AO221D0BWP7T port map(A1 => n_363, A2 => FE_OFN4_TL00_writeint, B1 => n_1, B2 => FE_PHN100_char2posx_3, C => n_12, Z => n_367);
  g7221 : MOAI22D0BWP7T port map(A1 => n_364, A2 => n_127, B1 => n_127, B2 => FE_PHN54_char1posxin_3, ZN => n_366);
  g7222 : ND2D1BWP7T port map(A1 => n_363, A2 => n_359, ZN => n_365);
  g7223 : INVD1BWP7T port map(I => n_364, ZN => n_363);
  g7224 : FA1D0BWP7T port map(A => n_322, B => n_52, CI => n_357, CO => n_362, S => n_364);
  g7227 : MOAI22D0BWP7T port map(A1 => n_359, A2 => n_59, B1 => n_61, B2 => FE_PHN85_char2posx_2, ZN => n_361);
  g7228 : MOAI22D0BWP7T port map(A1 => n_359, A2 => n_127, B1 => n_127, B2 => char1posxin(2), ZN => n_360);
  g7229 : INVD0BWP7T port map(I => n_359, ZN => n_358);
  g7230 : FA1D0BWP7T port map(A => n_319, B => n_50, CI => n_352, CO => n_357, S => n_359);
  g7233 : OAI211D1BWP7T port map(A1 => n_1, A2 => n_353, B => n_13, C => n_10, ZN => n_356);
  g7234 : MOAI22D0BWP7T port map(A1 => n_353, A2 => n_127, B1 => n_127, B2 => FE_PHN55_char1posxin_1, ZN => n_355);
  g7235 : NR2XD0BWP7T port map(A1 => n_353, A2 => n_328, ZN => n_354);
  g7236 : FA1D0BWP7T port map(A => n_321, B => n_55, CI => n_329, CO => n_352, S => n_353);
  g7245 : MOAI22D0BWP7T port map(A1 => n_328, A2 => n_127, B1 => n_127, B2 => char1posxin(0), ZN => n_351);
  g7246 : MOAI22D0BWP7T port map(A1 => n_328, A2 => n_59, B1 => n_61, B2 => FE_PHN164_char2posx_0, ZN => n_350);
  g7256 : MOAI22D0BWP7T port map(A1 => n_329, A2 => n_136, B1 => n_135, B2 => char1velxin(1), ZN => n_349);
  g7257 : MOAI22D0BWP7T port map(A1 => n_329, A2 => n_1, B1 => n_1, B2 => FE_PHN77_char2velx_1, ZN => n_348);
  g7262 : MOAI22D0BWP7T port map(A1 => n_317, A2 => n_1, B1 => n_1, B2 => FE_PHN75_char2velx_4, ZN => n_346);
  g7263 : MOAI22D0BWP7T port map(A1 => n_319, A2 => n_136, B1 => n_135, B2 => FE_PHN25_char1velxin_2, ZN => n_345);
  g7264 : AO22D0BWP7T port map(A1 => n_320, A2 => n_137, B1 => char1velxin(6), B2 => n_135, Z => n_344);
  g7265 : AO22D0BWP7T port map(A1 => n_324, A2 => n_137, B1 => FE_PHN61_char1velxin_8, B2 => n_135, Z => n_343);
  g7266 : MOAI22D0BWP7T port map(A1 => n_317, A2 => n_136, B1 => n_135, B2 => FE_PHN22_char1velxin_4, ZN => n_342);
  g7267 : MOAI22D0BWP7T port map(A1 => n_319, A2 => n_1, B1 => n_1, B2 => FE_PHN71_char2velx_2, ZN => n_341);
  g7269 : IND2D1BWP7T port map(A1 => n_331, B1 => n_330, ZN => n_347);
  g7270 : MOAI22D0BWP7T port map(A1 => n_323, A2 => n_1, B1 => n_1, B2 => FE_PHN66_char2velx_5, ZN => n_339);
  g7271 : MOAI22D0BWP7T port map(A1 => n_318, A2 => n_136, B1 => n_135, B2 => char1velxin(7), ZN => n_338);
  g7272 : MOAI22D0BWP7T port map(A1 => n_325, A2 => n_136, B1 => n_135, B2 => FE_PHN21_char1velxin_9, ZN => n_337);
  g7273 : MOAI22D0BWP7T port map(A1 => n_322, A2 => n_1, B1 => n_1, B2 => FE_PHN76_char2velx_3, ZN => n_336);
  g7274 : MOAI22D0BWP7T port map(A1 => n_323, A2 => n_136, B1 => n_135, B2 => FE_PHN27_char1velxin_5, ZN => n_335);
  g7275 : MOAI22D0BWP7T port map(A1 => n_318, A2 => n_1, B1 => n_1, B2 => FE_PHN70_char2velx_7, ZN => n_334);
  g7276 : MOAI22D0BWP7T port map(A1 => n_325, A2 => n_1, B1 => n_1, B2 => FE_PHN87_char2velx_9, ZN => n_333);
  g7277 : MOAI22D0BWP7T port map(A1 => n_322, A2 => n_136, B1 => n_135, B2 => char1velxin(3), ZN => n_332);
  g7278 : CKXOR2D1BWP7T port map(A1 => n_324, A2 => n_25, Z => n_340);
  g7279 : INR2D1BWP7T port map(A1 => n_320, B1 => n_39, ZN => n_331);
  g7280 : IND2D1BWP7T port map(A1 => n_320, B1 => n_39, ZN => n_330);
  g7281 : AOI21D0BWP7T port map(A1 => n_308, A2 => n_159, B => n_316, ZN => n_329);
  g7282 : MOAI22D0BWP7T port map(A1 => n_313, A2 => n_136, B1 => n_135, B2 => FE_PHN32_char1velxin_0, ZN => n_327);
  g7283 : MOAI22D0BWP7T port map(A1 => n_313, A2 => n_1, B1 => n_1, B2 => FE_PHN73_char2velx_0, ZN => n_326);
  g7284 : MAOI22D0BWP7T port map(A1 => n_312, A2 => n_63, B1 => n_312, B2 => n_63, ZN => n_328);
  g7285 : AOI21D0BWP7T port map(A1 => n_309, A2 => n_295, B => n_315, ZN => n_325);
  g7286 : IND2D1BWP7T port map(A1 => n_63, B1 => n_312, ZN => n_321);
  g7287 : OAI211D1BWP7T port map(A1 => n_505, A2 => n_306, B => n_314, C => n_310, ZN => n_324);
  g7288 : AOI221D0BWP7T port map(A1 => n_308, A2 => n_261, B1 => n_305, B2 => n_259, C => n_315, ZN => n_323);
  g7289 : AOI221D0BWP7T port map(A1 => n_308, A2 => n_201, B1 => n_305, B2 => n_197, C => n_315, ZN => n_322);
  g7290 : OAI22D0BWP7T port map(A1 => n_311, A2 => n_116, B1 => n_306, B2 => n_159, ZN => n_316);
  g7291 : OAI221D0BWP7T port map(A1 => n_307, A2 => n_273, B1 => n_271, B2 => n_306, C => n_314, ZN => n_320);
  g7292 : AOI221D0BWP7T port map(A1 => n_308, A2 => n_173, B1 => n_305, B2 => n_178, C => n_315, ZN => n_319);
  g7293 : AOI221D0BWP7T port map(A1 => n_308, A2 => n_279, B1 => n_305, B2 => n_284, C => n_315, ZN => n_318);
  g7294 : AOI221D0BWP7T port map(A1 => n_308, A2 => n_229, B1 => n_305, B2 => n_228, C => n_315, ZN => n_317);
  g7295 : INVD0BWP7T port map(I => n_315, ZN => n_314);
  g7296 : NR2D1BWP7T port map(A1 => n_311, A2 => n_79, ZN => n_315);
  g7297 : INVD0BWP7T port map(I => n_313, ZN => n_312);
  g7298 : OAI21D0BWP7T port map(A1 => n_308, A2 => n_305, B => n_122, ZN => n_313);
  g7299 : ND4D0BWP7T port map(A1 => n_303, A2 => n_302, A3 => n_206, A4 => n_122, ZN => n_311);
  g7300 : ND3D0BWP7T port map(A1 => n_308, A2 => n_292, A3 => n_278, ZN => n_310);
  g7301 : ND3D0BWP7T port map(A1 => n_307, A2 => n_292, A3 => n_285, ZN => n_309);
  g7302 : INVD0BWP7T port map(I => n_308, ZN => n_307);
  g7303 : OAI31D1BWP7T port map(A1 => n_281, A2 => n_283, A3 => n_300, B => n_304, ZN => n_308);
  g7304 : INVD1BWP7T port map(I => n_306, ZN => n_305);
  g7305 : OAI21D0BWP7T port map(A1 => n_300, A2 => n_288, B => n_304, ZN => n_306);
  g7306 : AOI31D0BWP7T port map(A1 => n_299, A2 => n_292, A3 => n_79, B => n_297, ZN => n_304);
  g7307 : AOI21D0BWP7T port map(A1 => n_301, A2 => n_288, B => n_298, ZN => n_303);
  g7308 : MAOI22D0BWP7T port map(A1 => n_199, A2 => n_151, B1 => n_301, B2 => n_288, ZN => n_302);
  g7309 : NR2D0BWP7T port map(A1 => n_296, A2 => n_297, ZN => n_301);
  g7310 : INVD0BWP7T port map(I => n_299, ZN => n_300);
  g7311 : AO221D0BWP7T port map(A1 => n_287, A2 => n_260, B1 => n_289, B2 => n_292, C => n_293, Z => n_298);
  g7312 : IAO21D0BWP7T port map(A1 => n_292, A2 => n_79, B => n_296, ZN => n_299);
  g7313 : NR2D1BWP7T port map(A1 => n_295, A2 => n_79, ZN => n_297);
  g7314 : AN2D0BWP7T port map(A1 => n_295, A2 => n_79, Z => n_296);
  g7315 : MOAI22D0BWP7T port map(A1 => n_290, A2 => n_120, B1 => n_290, B2 => n_120, ZN => n_295);
  g7317 : OAI22D0BWP7T port map(A1 => n_289, A2 => n_292, B1 => n_286, B2 => n_260, ZN => n_293);
  g7319 : FA1D0BWP7T port map(A => TL02_n_454, B => n_19, CI => n_274, CO => n_290, S => n_292);
  g7320 : OR2D1BWP7T port map(A1 => n_288, A2 => n_79, Z => n_289);
  g7321 : IAO21D0BWP7T port map(A1 => n_281, A2 => n_209, B => n_282, ZN => n_288);
  g7322 : ND4D0BWP7T port map(A1 => n_280, A2 => n_272, A3 => n_232, A4 => n_209, ZN => n_287);
  g7323 : NR4D0BWP7T port map(A1 => n_280, A2 => n_272, A3 => n_232, A4 => n_209, ZN => n_286);
  g7324 : HA1D0BWP7T port map(A => n_269, B => n_276, CO => n_285, S => n_284);
  g7325 : AOI211D0BWP7T port map(A1 => n_200, A2 => n_157, B => n_282, C => n_203, ZN => n_283);
  g7326 : NR2D1BWP7T port map(A1 => n_277, A2 => n_2, ZN => n_282);
  g7327 : AOI31D0BWP7T port map(A1 => n_276, A2 => n_268, A3 => n_256, B => n_79, ZN => n_281);
  g7328 : OAI21D0BWP7T port map(A1 => n_275, A2 => n_270, B => n_278, ZN => n_279);
  g7329 : MOAI22D0BWP7T port map(A1 => n_276, A2 => n_79, B1 => n_276, B2 => n_79, ZN => n_280);
  g7330 : ND2D1BWP7T port map(A1 => n_275, A2 => n_270, ZN => n_278);
  g7331 : NR4D0BWP7T port map(A1 => n_276, A2 => n_268, A3 => n_247, A4 => n_220, ZN => n_277);
  g7332 : INVD0BWP7T port map(I => n_276, ZN => n_275);
  g7333 : FA1D0BWP7T port map(A => TL02_n_456, B => n_53, CI => n_267, CO => n_274, S => n_276);
  g7334 : AOI21D0BWP7T port map(A1 => n_268, A2 => n_258, B => n_270, ZN => n_273);
  g7335 : MAOI22D0BWP7T port map(A1 => n_268, A2 => n_257, B1 => n_268, B2 => n_257, ZN => n_271);
  g7336 : MOAI22D0BWP7T port map(A1 => n_268, A2 => n_79, B1 => n_268, B2 => n_79, ZN => n_272);
  g7337 : NR2D1BWP7T port map(A1 => n_268, A2 => n_258, ZN => n_270);
  g7338 : INR2XD0BWP7T port map(A1 => n_268, B1 => n_257, ZN => n_269);
  g7339 : FA1D0BWP7T port map(A => TL02_n_457, B => n_18, CI => n_244, CO => n_267, S => n_268);
  g7342 : AO22D0BWP7T port map(A1 => n_262, A2 => n_137, B1 => FE_PHN46_char1posyin_7, B2 => n_135, Z => n_266);
  g7343 : AO22D0BWP7T port map(A1 => n_262, A2 => n_60, B1 => FE_PHN168_char2posy_7, B2 => n_61, Z => n_265);
  g7344 : ND3D0BWP7T port map(A1 => n_251, A2 => n_238, A3 => n_183, ZN => n_264);
  g7345 : OAI211D1BWP7T port map(A1 => n_245, A2 => n_250, B => n_249, C => n_253, ZN => n_263);
  g7346 : OAI21D0BWP7T port map(A1 => n_246, A2 => n_222, B => n_258, ZN => n_261);
  g7347 : IND2D1BWP7T port map(A1 => n_243, B1 => n_252, ZN => n_262);
  g7348 : MOAI22D0BWP7T port map(A1 => n_247, A2 => n_223, B1 => n_247, B2 => n_223, ZN => n_259);
  g7349 : OAI22D0BWP7T port map(A1 => n_247, A2 => n_79, B1 => n_246, B2 => n_2, ZN => n_260);
  g7350 : INR2D0BWP7T port map(A1 => n_220, B1 => n_246, ZN => n_256);
  g7351 : IAO21D0BWP7T port map(A1 => n_183, A2 => n_166, B => n_245, ZN => n_255);
  g7352 : OAI31D0BWP7T port map(A1 => n_207, A2 => n_215, A3 => n_231, B => n_243, ZN => n_254);
  g7353 : ND2D1BWP7T port map(A1 => n_246, A2 => n_222, ZN => n_258);
  g7354 : IND2D1BWP7T port map(A1 => n_223, B1 => n_247, ZN => n_257);
  g7355 : CKND1BWP7T port map(I => n_251, ZN => n_250);
  g7356 : AOI222D0BWP7T port map(A1 => n_239, A2 => n_164, B1 => inputsp1(3), B2 => FE_OFN0_n_6, C1 => inputsp2(3), C2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_249);
  g7357 : AOI211XD0BWP7T port map(A1 => n_162, A2 => n_139, B => n_242, C => n_208, ZN => n_248);
  g7358 : MAOI22D0BWP7T port map(A1 => n_235, A2 => n_142, B1 => n_235, B2 => n_142, ZN => n_253);
  g7359 : MAOI22D0BWP7T port map(A1 => n_240, A2 => n_237, B1 => n_240, B2 => n_237, ZN => n_252);
  g7360 : MOAI22D0BWP7T port map(A1 => n_231, A2 => n_233, B1 => n_231, B2 => n_233, ZN => n_251);
  g7361 : INVD1BWP7T port map(I => n_247, ZN => n_246);
  g7362 : FA1D0BWP7T port map(A => TL02_n_458, B => n_17, CI => n_217, CO => n_244, S => n_247);
  g7363 : ND2D1BWP7T port map(A1 => n_238, A2 => n_213, ZN => n_245);
  g7364 : MOAI22D0BWP7T port map(A1 => n_234, A2 => n_241, B1 => n_234, B2 => n_241, ZN => n_243);
  g7365 : INVD0BWP7T port map(I => n_238, ZN => n_242);
  g7366 : AN4D0BWP7T port map(A1 => n_216, A2 => n_205, A3 => n_184, A4 => n_147, Z => n_239);
  g7367 : AOI21D0BWP7T port map(A1 => n_211, A2 => n_224, B => n_210, ZN => n_241);
  g7368 : AO21D0BWP7T port map(A1 => n_225, A2 => n_226, B => n_227, Z => n_240);
  g7369 : MOAI22D0BWP7T port map(A1 => n_214, A2 => n_208, B1 => n_214, B2 => n_208, ZN => n_238);
  g7370 : MAOI22D0BWP7T port map(A1 => n_221, A2 => n_125, B1 => n_221, B2 => n_125, ZN => n_237);
  g7371 : MAOI22D0BWP7T port map(A1 => n_219, A2 => n_224, B1 => n_219, B2 => n_224, ZN => n_236);
  g7372 : INR2XD0BWP7T port map(A1 => n_221, B1 => n_125, ZN => n_235);
  g7373 : INR2D1BWP7T port map(A1 => n_226, B1 => n_227, ZN => n_234);
  g7374 : ND2D1BWP7T port map(A1 => n_215, A2 => n_208, ZN => n_233);
  g7375 : INVD0BWP7T port map(I => n_231, ZN => n_230);
  g7376 : AO21D0BWP7T port map(A1 => n_220, A2 => n_196, B => n_222, Z => n_229);
  g7377 : MOAI22D0BWP7T port map(A1 => n_220, A2 => n_194, B1 => n_220, B2 => n_194, ZN => n_228);
  g7378 : MOAI22D0BWP7T port map(A1 => n_220, A2 => n_79, B1 => n_220, B2 => n_79, ZN => n_232);
  g7379 : MOAI22D0BWP7T port map(A1 => n_218, A2 => n_191, B1 => n_218, B2 => n_191, ZN => n_231);
  g7380 : AO21D0BWP7T port map(A1 => n_211, A2 => n_202, B => n_210, Z => n_225);
  g7381 : NR2XD0BWP7T port map(A1 => n_216, A2 => n_46, ZN => n_227);
  g7382 : ND2D1BWP7T port map(A1 => n_216, A2 => n_46, ZN => n_226);
  g7383 : OAI21D0BWP7T port map(A1 => n_212, A2 => n_185, B => n_195, ZN => n_224);
  g7384 : IND2D1BWP7T port map(A1 => n_194, B1 => n_220, ZN => n_223);
  g7385 : NR2D1BWP7T port map(A1 => n_220, A2 => n_196, ZN => n_222);
  g7386 : OAI211D1BWP7T port map(A1 => n_133, A2 => n_204, B => n_132, C => n_87, ZN => n_221);
  g7387 : FA1D0BWP7T port map(A => TL02_n_459, B => n_20, CI => n_190, CO => n_217, S => n_220);
  g7388 : IND2D1BWP7T port map(A1 => n_210, B1 => n_211, ZN => n_219);
  g7389 : IND2D1BWP7T port map(A1 => n_176, B1 => n_212, ZN => n_218);
  g7390 : INVD1BWP7T port map(I => n_215, ZN => n_214);
  g7391 : OAI21D0BWP7T port map(A1 => n_198, A2 => n_183, B => n_208, ZN => n_213);
  g7392 : MAOI22D0BWP7T port map(A1 => n_204, A2 => n_144, B1 => n_204, B2 => n_144, ZN => n_216);
  g7393 : MOAI22D0BWP7T port map(A1 => n_177, A2 => n_188, B1 => n_177, B2 => n_188, ZN => n_215);
  g7394 : ND2D1BWP7T port map(A1 => n_175, A2 => n_188, ZN => n_212);
  g7395 : ND2D1BWP7T port map(A1 => n_205, A2 => n_44, ZN => n_211);
  g7396 : NR2XD0BWP7T port map(A1 => n_205, A2 => n_44, ZN => n_210);
  g7397 : IAO21D0BWP7T port map(A1 => n_182, A2 => n_166, B => n_198, ZN => n_207);
  g7398 : CKMUX2D1BWP7T port map(I0 => n_199, I1 => n_151, S => n_172, Z => n_206);
  g7399 : AOI21D0BWP7T port map(A1 => n_200, A2 => n_150, B => n_203, ZN => n_209);
  g7400 : ND2D1BWP7T port map(A1 => n_198, A2 => n_183, ZN => n_208);
  g7401 : FA1D0BWP7T port map(A => n_121, B => n_84, CI => n_171, CO => n_204, S => n_205);
  g7402 : IND2D1BWP7T port map(A1 => n_175, B1 => n_195, ZN => n_202);
  g7403 : OAI21D0BWP7T port map(A1 => n_193, A2 => n_170, B => n_196, ZN => n_201);
  g7404 : AOI21D0BWP7T port map(A1 => n_193, A2 => n_163, B => n_2, ZN => n_203);
  g7405 : MOAI22D0BWP7T port map(A1 => n_193, A2 => n_179, B1 => n_193, B2 => n_179, ZN => n_197);
  g7406 : OAI21D0BWP7T port map(A1 => n_193, A2 => n_163, B => n_2, ZN => n_200);
  g7407 : MAOI22D0BWP7T port map(A1 => n_193, A2 => n_2, B1 => n_193, B2 => n_2, ZN => n_199);
  g7408 : MAOI22D0BWP7T port map(A1 => n_506, A2 => n_164, B1 => n_506, B2 => n_164, ZN => n_198);
  g7409 : ND2D1BWP7T port map(A1 => n_193, A2 => n_170, ZN => n_196);
  g7410 : AOI21D0BWP7T port map(A1 => n_186, A2 => n_176, B => n_187, ZN => n_195);
  g7411 : ND2D1BWP7T port map(A1 => n_192, A2 => n_179, ZN => n_194);
  g7412 : INVD1BWP7T port map(I => n_192, ZN => n_193);
  g7413 : FA1D0BWP7T port map(A => TL02_n_460, B => n_21, CI => n_154, CO => n_190, S => n_192);
  g7414 : IND2D1BWP7T port map(A1 => n_187, B1 => n_186, ZN => n_191);
  g7416 : MAOI222D1BWP7T port map(A => n_180, B => n_164, C => n_34, ZN => n_188);
  g7417 : NR2D1BWP7T port map(A1 => n_174, A2 => n_41, ZN => n_187);
  g7418 : INVD0BWP7T port map(I => n_186, ZN => n_185);
  g7419 : AN4D0BWP7T port map(A1 => n_174, A2 => n_169, A3 => n_138, A4 => n_115, Z => n_184);
  g7420 : ND2D1BWP7T port map(A1 => n_174, A2 => n_41, ZN => n_186);
  g7421 : INVD0BWP7T port map(I => n_183, ZN => n_182);
  g7423 : FA1D0BWP7T port map(A => n_161, B => n_22, CI => n_147, CO => n_180, S => n_183);
  g7424 : HA1D0BWP7T port map(A => n_153, B => n_168, CO => n_179, S => n_178);
  g7425 : IND2D1BWP7T port map(A1 => n_176, B1 => n_175, ZN => n_177);
  g7426 : NR2XD0BWP7T port map(A1 => n_169, A2 => n_40, ZN => n_176);
  g7427 : ND2D1BWP7T port map(A1 => n_169, A2 => n_40, ZN => n_175);
  g7428 : AO21D0BWP7T port map(A1 => n_168, A2 => n_152, B => n_170, Z => n_173);
  g7429 : OAI22D0BWP7T port map(A1 => n_168, A2 => n_79, B1 => n_163, B2 => n_2, ZN => n_172);
  g7430 : MAOI22D0BWP7T port map(A1 => n_167, A2 => n_124, B1 => n_167, B2 => n_124, ZN => n_174);
  g7431 : IND2D1BWP7T port map(A1 => n_124, B1 => n_167, ZN => n_171);
  g7432 : NR2D1BWP7T port map(A1 => n_168, A2 => n_152, ZN => n_170);
  g7433 : MAOI22D0BWP7T port map(A1 => n_165, A2 => n_83, B1 => n_165, B2 => n_83, ZN => n_169);
  g7434 : INVD1BWP7T port map(I => n_163, ZN => n_168);
  g7435 : MOAI22D0BWP7T port map(A1 => n_160, A2 => n_117, B1 => TL02_n_597, B2 => n_36, ZN => n_167);
  g7436 : NR2D1BWP7T port map(A1 => n_162, A2 => n_139, ZN => n_166);
  g7437 : MOAI22D0BWP7T port map(A1 => n_158, A2 => n_117, B1 => n_158, B2 => n_117, ZN => n_165);
  g7438 : MAOI22D0BWP7T port map(A1 => n_156, A2 => n_81, B1 => n_156, B2 => n_81, ZN => n_164);
  g7439 : MAOI22D0BWP7T port map(A1 => n_507, A2 => TL02_n_461, B1 => n_507, B2 => TL02_n_461, ZN => n_163);
  g7440 : FA1D0BWP7T port map(A => n_134, B => n_24, CI => n_138, CO => n_161, S => n_162);
  g7441 : INR2D1BWP7T port map(A1 => n_158, B1 => n_83, ZN => n_160);
  g7442 : IOA21D0BWP7T port map(A1 => n_146, A2 => n_116, B => n_122, ZN => n_157);
  g7443 : IND2D1BWP7T port map(A1 => n_153, B1 => n_152, ZN => n_159);
  g7444 : OAI21D0BWP7T port map(A1 => n_148, A2 => n_81, B => n_123, ZN => n_158);
  g7445 : MOAI22D0BWP7T port map(A1 => n_148, A2 => n_123, B1 => n_148, B2 => n_123, ZN => n_156);
  g7447 : MAOI222D1BWP7T port map(A => n_140, B => n_4, C => n_31, ZN => n_154);
  g7448 : INR2XD0BWP7T port map(A1 => n_146, B1 => n_122, ZN => n_153);
  g7449 : INVD1BWP7T port map(I => n_151, ZN => n_150);
  g7450 : IND2D1BWP7T port map(A1 => n_146, B1 => n_122, ZN => n_152);
  g7451 : NR2XD0BWP7T port map(A1 => n_146, A2 => n_116, ZN => n_151);
  g7453 : OAI21D0BWP7T port map(A1 => n_131, A2 => n_130, B => n_143, ZN => n_148);
  g7454 : MAOI22D0BWP7T port map(A1 => n_145, A2 => n_130, B1 => n_145, B2 => n_130, ZN => n_147);
  g7455 : MOAI22D0BWP7T port map(A1 => n_141, A2 => TL02_n_462, B1 => n_141, B2 => TL02_n_462, ZN => n_146);
  g7456 : INR2XD0BWP7T port map(A1 => n_143, B1 => n_131, ZN => n_145);
  g7457 : INR2XD0BWP7T port map(A1 => n_132, B1 => n_133, ZN => n_144);
  g7458 : IND3D1BWP7T port map(A1 => n_81, B1 => n_128, B2 => n_86, ZN => n_143);
  g7459 : MOAI22D0BWP7T port map(A1 => n_118, A2 => n_76, B1 => n_118, B2 => n_76, ZN => n_142);
  g7460 : MAOI22D0BWP7T port map(A1 => n_82, A2 => n_33, B1 => n_82, B2 => n_33, ZN => n_141);
  g7461 : MAOI222D1BWP7T port map(A => TL02_n_462, B => n_82, C => n_32, ZN => n_140);
  g7462 : XNR2D1BWP7T port map(A1 => n_115, A2 => n_38, ZN => n_139);
  g7463 : MAOI22D0BWP7T port map(A1 => n_129, A2 => n_77, B1 => n_129, B2 => n_77, ZN => n_138);
  g7464 : INVD1BWP7T port map(I => n_137, ZN => n_136);
  g7465 : OR2D1BWP7T port map(A1 => n_115, A2 => n_38, Z => n_134);
  g7466 : NR2XD0BWP7T port map(A1 => n_127, A2 => FE_OFN3_reset, ZN => n_137);
  g7467 : NR2D1P5BWP7T port map(A1 => n_126, A2 => FE_OFN3_reset, ZN => n_135);
  g7468 : NR2D1BWP7T port map(A1 => n_85, A2 => n_119, ZN => n_133);
  g7469 : ND2D1BWP7T port map(A1 => n_85, A2 => n_119, ZN => n_132);
  g7470 : AOI21D0BWP7T port map(A1 => n_86, A2 => n_80, B => n_128, ZN => n_131);
  g7471 : IND2D1BWP7T port map(A1 => n_77, B1 => n_129, ZN => n_130);
  g7473 : HA1D0BWP7T port map(A => n_23, B => TL02_n_600, CO => n_128, S => n_129);
  g7488 : INVD0BWP7T port map(I => n_127, ZN => n_126);
  g7502 : ND4D1BWP7T port map(A1 => n_68, A2 => n_29, A3 => n_28, A4 => n_26, ZN => n_127);
  g7504 : AO21D0BWP7T port map(A1 => n_5, A2 => n_45, B => n_85, Z => n_121);
  g7525 : AO21D0BWP7T port map(A1 => n_3, A2 => n_65, B => n_76, Z => n_125);
  g7531 : OAI21D0BWP7T port map(A1 => TL02_n_596, A2 => n_47, B => n_84, ZN => n_124);
  g7532 : IAO21D0BWP7T port map(A1 => TL02_n_598, A2 => n_43, B => n_83, ZN => n_123);
  g7534 : AO21D0BWP7T port map(A1 => n_9, A2 => n_64, B => n_82, Z => n_122);
  g7536 : AO22D0BWP7T port map(A1 => n_57, A2 => char1perc(4), B1 => n_58, B2 => char1percin(4), Z => n_114);
  g7537 : AO22D0BWP7T port map(A1 => n_57, A2 => char1posx(4), B1 => FE_PHN50_char1posxin_4, B2 => n_58, Z => n_113);
  g7538 : AO22D0BWP7T port map(A1 => n_57, A2 => char1posx(8), B1 => FE_PHN52_char1posxin_8, B2 => n_58, Z => n_112);
  g7539 : AO22D0BWP7T port map(A1 => n_57, A2 => char1posy(0), B1 => char1posyin(0), B2 => n_58, Z => n_111);
  g7540 : AO22D0BWP7T port map(A1 => n_57, A2 => FE_PHN110_char1perc_0, B1 => char1percin(0), B2 => n_58, Z => n_110);
  g7541 : AO22D0BWP7T port map(A1 => n_57, A2 => char1posx(7), B1 => char1posxin(7), B2 => n_58, Z => n_109);
  g7542 : AO22D0BWP7T port map(A1 => n_57, A2 => char1posy(1), B1 => char1posyin(1), B2 => n_58, Z => n_108);
  g7543 : AO22D0BWP7T port map(A1 => n_57, A2 => char1posy(3), B1 => char1posyin(3), B2 => n_58, Z => FE_PHN136_n_107);
  g7544 : AO22D0BWP7T port map(A1 => n_61, A2 => FE_PHN118_char2perc_1, B1 => n_60, B2 => char2percin(1), Z => n_106);
  g7545 : AO22D0BWP7T port map(A1 => n_57, A2 => char1posy(4), B1 => char1posyin(4), B2 => n_58, Z => n_105);
  g7546 : AO22D0BWP7T port map(A1 => n_61, A2 => char2perc(4), B1 => n_60, B2 => char2percin(4), Z => n_104);
  g7547 : AO22D0BWP7T port map(A1 => n_61, A2 => FE_PHN90_char2perc_3, B1 => n_60, B2 => char2percin(3), Z => n_103);
  g7548 : AO22D0BWP7T port map(A1 => n_57, A2 => char1perc(1), B1 => n_58, B2 => char1percin(1), Z => n_102);
  g7549 : AO22D0BWP7T port map(A1 => n_57, A2 => char1posx(5), B1 => FE_PHN69_char1posxin_5, B2 => n_58, Z => FE_PHN140_n_101);
  g7550 : AO22D0BWP7T port map(A1 => n_57, A2 => char1perc(2), B1 => n_58, B2 => char1percin(2), Z => n_100);
  g7551 : AO22D0BWP7T port map(A1 => n_57, A2 => char1posy(7), B1 => FE_PHN46_char1posyin_7, B2 => n_58, Z => n_99);
  g7552 : AO22D0BWP7T port map(A1 => n_57, A2 => char1posx(3), B1 => FE_PHN54_char1posxin_3, B2 => n_58, Z => n_98);
  g7553 : AO22D0BWP7T port map(A1 => n_57, A2 => char1perc(3), B1 => n_58, B2 => char1percin(3), Z => n_97);
  g7554 : AO22D0BWP7T port map(A1 => n_57, A2 => char1perc(5), B1 => n_58, B2 => char1percin(5), Z => n_96);
  g7555 : AO22D0BWP7T port map(A1 => n_57, A2 => char1perc(6), B1 => n_58, B2 => char1percin(6), Z => n_95);
  g7556 : AO22D0BWP7T port map(A1 => n_57, A2 => FE_PHN112_char1perc_7, B1 => n_58, B2 => char1percin(7), Z => n_94);
  g7557 : AO22D0BWP7T port map(A1 => n_61, A2 => FE_PHN102_char2perc_0, B1 => char2percin(0), B2 => n_60, Z => n_93);
  g7558 : AO22D0BWP7T port map(A1 => n_61, A2 => FE_PHN97_char2perc_2, B1 => n_60, B2 => char2percin(2), Z => n_92);
  g7559 : AO22D0BWP7T port map(A1 => n_61, A2 => char2perc(5), B1 => n_60, B2 => char2percin(5), Z => n_91);
  g7560 : AO22D0BWP7T port map(A1 => n_61, A2 => char2perc(6), B1 => n_60, B2 => char2percin(6), Z => n_90);
  g7561 : AO22D0BWP7T port map(A1 => n_61, A2 => FE_PHN117_char2perc_7, B1 => n_60, B2 => char2percin(7), Z => n_89);
  g7562 : AO22D0BWP7T port map(A1 => n_57, A2 => char1posx(0), B1 => char1posxin(0), B2 => n_58, Z => n_88);
  g7563 : CKXOR2D1BWP7T port map(A1 => TL02_n_454, A2 => n_54, Z => n_120);
  g7564 : OA21D0BWP7T port map(A1 => TL02_n_594, A2 => n_67, B => n_87, Z => n_119);
  g7565 : MOAI22D0BWP7T port map(A1 => TL02_n_592, A2 => n_48, B1 => TL02_n_592, B2 => n_48, ZN => n_118);
  g7566 : MAOI22D0BWP7T port map(A1 => TL02_n_597, A2 => n_35, B1 => TL02_n_597, B2 => n_35, ZN => n_117);
  g7567 : AOI21D0BWP7T port map(A1 => n_49, A2 => n_66, B => n_2, ZN => n_116);
  g7568 : MOAI22D0BWP7T port map(A1 => TL02_n_601, A2 => n_37, B1 => TL02_n_601, B2 => n_37, ZN => n_115);
  g7569 : INVD1BWP7T port map(I => n_80, ZN => n_81);
  g7570 : INVD1BWP7T port map(I => n_2, ZN => n_79);
  g7571 : ND2D0BWP7T port map(A1 => n_61, A2 => FE_PHN95_char2posy_0, ZN => n_78);
  g7572 : ND2D1BWP7T port map(A1 => TL02_n_594, A2 => n_67, ZN => n_87);
  g7573 : IND2D1BWP7T port map(A1 => TL02_n_599, B1 => n_42, ZN => n_86);
  g7574 : NR2XD0BWP7T port map(A1 => n_5, A2 => n_45, ZN => n_85);
  g7575 : ND2D1BWP7T port map(A1 => TL02_n_596, A2 => n_47, ZN => n_84);
  g7576 : AN2D1BWP7T port map(A1 => TL02_n_598, A2 => n_43, Z => n_83);
  g7577 : NR2D1BWP7T port map(A1 => n_9, A2 => n_64, ZN => n_82);
  g7578 : IND2D1BWP7T port map(A1 => n_42, B1 => TL02_n_599, ZN => n_80);
  g7579 : NR2XD0BWP7T port map(A1 => n_49, A2 => n_66, ZN => n_2);
  g7580 : AO221D0BWP7T port map(A1 => n_1, A2 => char1posx(1), B1 => FE_OFN4_TL00_writeint, B2 => FE_PHN55_char1posxin_1, C => n_15, Z => n_75);
  g7581 : AO221D0BWP7T port map(A1 => n_1, A2 => char1posy(5), B1 => FE_OFN4_TL00_writeint, B2 => char1posyin(5), C => n_15, Z => n_74);
  g7582 : AO221D0BWP7T port map(A1 => n_1, A2 => char1posy(6), B1 => FE_OFN4_TL00_writeint, B2 => char1posyin(6), C => n_15, Z => FE_PHN143_n_73);
  g7583 : AO221D0BWP7T port map(A1 => n_1, A2 => char1posx(2), B1 => FE_OFN4_TL00_writeint, B2 => char1posxin(2), C => n_15, Z => n_72);
  g7584 : AO221D0BWP7T port map(A1 => n_1, A2 => char1posy(2), B1 => FE_OFN4_TL00_writeint, B2 => char1posyin(2), C => n_15, Z => FE_PHN138_n_71);
  g7585 : AO221D0BWP7T port map(A1 => n_1, A2 => char1posx(6), B1 => FE_OFN4_TL00_writeint, B2 => FE_PHN67_char1posxin_6, C => n_15, Z => n_70);
  g7586 : NR4D0BWP7T port map(A1 => FE_OFN4_TL00_writeint, A2 => FE_PHN58_TL00_WL00_state_1, A3 => Vsync, A4 => FE_OFN3_reset, ZN => n_69);
  g7587 : IINR4D0BWP7T port map(A1 => n_508, A2 => vcountintern(8), B1 => vcountintern(9), B2 => hcountintern(1), ZN => n_68);
  g7588 : INR2XD0BWP7T port map(A1 => n_37, B1 => TL02_n_601, ZN => n_77);
  g7589 : NR2XD0BWP7T port map(A1 => n_3, A2 => n_65, ZN => n_76);
  g7590 : INVD1BWP7T port map(I => n_60, ZN => n_59);
  g7605 : IOA21D0BWP7T port map(A1 => FE_PHN58_TL00_WL00_state_1, A2 => TL01_n_63, B => n_1, ZN => n_56);
  g7606 : AOI22D0BWP7T port map(A1 => char1posx(1), A2 => FE_OFN0_n_6, B1 => char2posx(1), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_55);
  g7607 : OAI22D0BWP7T port map(A1 => char1velx(9), A2 => FE_OFN1_TL02_PHS0_sel_0, B1 => FE_PHN176_char2velx_9, B2 => FE_OFN0_n_6, ZN => n_54);
  g7608 : OA22D0BWP7T port map(A1 => char1vely(7), A2 => FE_OFN1_TL02_PHS0_sel_0, B1 => FE_OFN0_n_6, B2 => char2vely(7), Z => n_67);
  g7609 : AO22D0BWP7T port map(A1 => inputsp1(1), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => inputsp2(1), Z => n_66);
  g7610 : AOI22D0BWP7T port map(A1 => char1vely(8), A2 => FE_OFN0_n_6, B1 => char2vely(8), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_65);
  g7611 : OAI22D0BWP7T port map(A1 => char1velx(0), A2 => FE_OFN1_TL02_PHS0_sel_0, B1 => char2velx(0), B2 => FE_OFN0_n_6, ZN => n_64);
  g7612 : AOI22D0BWP7T port map(A1 => char1posx(0), A2 => FE_OFN0_n_6, B1 => char2posx(0), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_63);
  g7613 : AO22D0BWP7T port map(A1 => char1velx(7), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => char2velx(7), Z => n_53);
  g7614 : AOI22D0BWP7T port map(A1 => char1posx(3), A2 => FE_OFN0_n_6, B1 => char2posx(3), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_52);
  g7615 : AOI22D0BWP7T port map(A1 => char1posx(5), A2 => FE_OFN0_n_6, B1 => char2posx(5), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_62);
  g7616 : AOI22D0BWP7T port map(A1 => char1posx(4), A2 => FE_OFN0_n_6, B1 => char2posx(4), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_51);
  g7617 : AOI22D0BWP7T port map(A1 => char1posx(2), A2 => FE_OFN0_n_6, B1 => char2posx(2), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_50);
  g7618 : NR2XD0BWP7T port map(A1 => n_12, A2 => FE_OFN4_TL00_writeint, ZN => n_61);
  g7619 : NR2XD0BWP7T port map(A1 => n_12, A2 => n_1, ZN => n_60);
  g7620 : NR2XD0BWP7T port map(A1 => n_15, A2 => n_1, ZN => n_58);
  g7621 : NR2XD0BWP7T port map(A1 => n_15, A2 => FE_OFN4_TL00_writeint, ZN => n_57);
  g7622 : INVD0BWP7T port map(I => n_35, ZN => n_36);
  g7623 : INVD0BWP7T port map(I => n_33, ZN => n_32);
  g7624 : IINR4D0BWP7T port map(A1 => vcountintern(1), A2 => vcountintern(2), B1 => vcountintern(3), B2 => vcountintern(0), ZN => n_29);
  g7625 : NR4D0BWP7T port map(A1 => hcountintern(8), A2 => hcountintern(9), A3 => hcountintern(7), A4 => hcountintern(6), ZN => n_28);
  g7627 : NR4D0BWP7T port map(A1 => hcountintern(5), A2 => hcountintern(4), A3 => hcountintern(3), A4 => hcountintern(2), ZN => n_26);
  g7628 : AOI22D0BWP7T port map(A1 => inputsp1(0), A2 => FE_OFN0_n_6, B1 => inputsp2(0), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_49);
  g7629 : OAI22D0BWP7T port map(A1 => char1posx(8), A2 => FE_OFN1_TL02_PHS0_sel_0, B1 => FE_PHN123_char2posx_8, B2 => FE_OFN0_n_6, ZN => n_25);
  g7630 : AOI22D0BWP7T port map(A1 => char1vely(9), A2 => FE_OFN0_n_6, B1 => char2vely(9), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_48);
  g7631 : OA22D0BWP7T port map(A1 => char1vely(5), A2 => FE_OFN1_TL02_PHS0_sel_0, B1 => FE_OFN0_n_6, B2 => char2vely(5), Z => n_47);
  g7632 : AOI22D0BWP7T port map(A1 => char1posy(7), A2 => FE_OFN0_n_6, B1 => char2posy(7), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_46);
  g7633 : OAI22D0BWP7T port map(A1 => char1vely(6), A2 => FE_OFN1_TL02_PHS0_sel_0, B1 => char2vely(6), B2 => FE_OFN0_n_6, ZN => n_45);
  g7634 : OAI22D0BWP7T port map(A1 => char1posy(6), A2 => FE_OFN1_TL02_PHS0_sel_0, B1 => char2posy(6), B2 => FE_OFN0_n_6, ZN => n_44);
  g7635 : AOI22D0BWP7T port map(A1 => char1posy(1), A2 => FE_OFN0_n_6, B1 => char2posy(1), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_24);
  g7636 : OA22D0BWP7T port map(A1 => char1vely(3), A2 => FE_OFN1_TL02_PHS0_sel_0, B1 => FE_OFN0_n_6, B2 => char2vely(3), Z => n_43);
  g7637 : AOI22D0BWP7T port map(A1 => char1vely(2), A2 => FE_OFN0_n_6, B1 => char2vely(2), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_42);
  g7638 : AOI22D0BWP7T port map(A1 => char1posy(5), A2 => FE_OFN0_n_6, B1 => char2posy(5), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_41);
  g7639 : OAI22D0BWP7T port map(A1 => char1posy(4), A2 => FE_OFN1_TL02_PHS0_sel_0, B1 => char2posy(4), B2 => FE_OFN0_n_6, ZN => n_40);
  g7640 : AOI22D0BWP7T port map(A1 => char1posx(6), A2 => FE_OFN0_n_6, B1 => char2posx(6), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_39);
  g7641 : AOI22D0BWP7T port map(A1 => char1posy(0), A2 => FE_OFN0_n_6, B1 => char2posy(0), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_38);
  g7642 : AOI22D0BWP7T port map(A1 => char1vely(0), A2 => FE_OFN0_n_6, B1 => char2vely(0), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_37);
  g7643 : AO22D0BWP7T port map(A1 => char1vely(1), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => char2vely(1), Z => n_23);
  g7644 : OAI22D0BWP7T port map(A1 => char1vely(4), A2 => FE_OFN1_TL02_PHS0_sel_0, B1 => char2vely(4), B2 => FE_OFN0_n_6, ZN => n_35);
  g7645 : AOI22D0BWP7T port map(A1 => char1posy(3), A2 => FE_OFN0_n_6, B1 => char2posy(3), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_34);
  g7646 : AOI22D0BWP7T port map(A1 => char1posy(2), A2 => FE_OFN0_n_6, B1 => char2posy(2), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_22);
  g7647 : AOI22D0BWP7T port map(A1 => char1velx(1), A2 => FE_OFN0_n_6, B1 => char2velx(1), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_33);
  g7648 : AO22D0BWP7T port map(A1 => char1velx(3), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => char2velx(3), Z => n_21);
  g7649 : AOI22D0BWP7T port map(A1 => char1velx(2), A2 => FE_OFN0_n_6, B1 => char2velx(2), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_31);
  g7650 : AO22D0BWP7T port map(A1 => char1velx(4), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => char2velx(4), Z => n_20);
  g7651 : AO22D0BWP7T port map(A1 => char1velx(8), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => char2velx(8), Z => n_19);
  g7652 : AOI22D0BWP7T port map(A1 => char1posx(7), A2 => FE_OFN0_n_6, B1 => char2posx(7), B2 => FE_OFN1_TL02_PHS0_sel_0, ZN => n_30);
  g7653 : AO22D0BWP7T port map(A1 => char1velx(6), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => char2velx(6), Z => n_18);
  g7654 : AO22D0BWP7T port map(A1 => char1velx(5), A2 => FE_OFN0_n_6, B1 => FE_OFN1_TL02_PHS0_sel_0, B2 => char2velx(5), Z => n_17);
  g7655 : INVD1BWP7T port map(I => n_16, ZN => n_15);
  g7656 : ND2D1BWP7T port map(A1 => n_1, A2 => FE_PHN82_char2posx_4, ZN => n_14);
  g7657 : NR2D1P5BWP7T port map(A1 => char1death, A2 => FE_OFN3_reset, ZN => n_16);
  g7658 : INVD1BWP7T port map(I => n_13, ZN => n_12);
  g7659 : ND2D1BWP7T port map(A1 => n_1, A2 => FE_PHN86_char2vely_3, ZN => n_11);
  g7660 : ND2D1BWP7T port map(A1 => n_1, A2 => FE_PHN165_char2posx_1, ZN => n_10);
  g7661 : NR2D1P5BWP7T port map(A1 => char2death, A2 => FE_OFN3_reset, ZN => n_13);
  g7662 : CKND1BWP7T port map(I => TL02_n_463, ZN => n_9);
  g7666 : INVD0BWP7T port map(I => TL02_n_595, ZN => n_5);
  g7667 : INVD0BWP7T port map(I => TL02_n_461, ZN => n_4);
  g7668 : INVD1BWP7T port map(I => TL02_n_592, ZN => n_3);
  TL00_WL00_state_reg_0 : DFD1BWP7T port map(CP => CTS_15, D => n_69, Q => TL00_writeint, QN => n_1);
  g2 : IND2D1BWP7T port map(A1 => n_432, B1 => n_137, ZN => n_0);
  g7672 : CKXOR2D1BWP7T port map(A1 => n_383, A2 => n_318, Z => n_504);
  g7673 : XNR2D1BWP7T port map(A1 => n_292, A2 => n_285, ZN => n_505);
  g7674 : CKXOR2D1BWP7T port map(A1 => n_180, A2 => n_34, Z => n_506);
  g7675 : XNR2D1BWP7T port map(A1 => n_140, A2 => n_31, ZN => n_507);
  g7676 : NR4D0BWP7T port map(A1 => vcountintern(6), A2 => vcountintern(7), A3 => vcountintern(5), A4 => vcountintern(4), ZN => n_508);
  TL02_PHS0_sel_reg_0 : DFD1BWP7T port map(CP => CTS_17, D => n_480, Q => TL02_PHS0_sel_0, QN => n_6);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1690 : OAI31D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_97, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_122, A3 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_171, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_173, ZN => TL02_n_592);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1691 : AO31D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_171, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_122, A3 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_97, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_96, Z => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_173);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1692 : MOAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_171, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_129, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_171, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_129, ZN => TL02_n_594);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1693 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_136, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_121, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_168, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_171, S => TL02_n_595);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1694 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_141, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_137, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_166, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_168, S => TL02_n_596);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1695 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_142, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_148, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_164, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_166, S => TL02_n_597);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1696 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_149, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_156, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_162, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_164, S => TL02_n_598);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1697 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_157, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_153, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_160, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_162, S => TL02_n_599);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1698 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_154, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_151, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_158, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_160, S => TL02_n_600);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1699 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_152, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_144, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_155, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_158, S => TL02_n_601);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1700 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_146, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_105, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_124, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_156, S => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_157);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1701 : MAOI222D1BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_150, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_143, C => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_134, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_155);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1702 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_138, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_109, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_147, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_153, S => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_154);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1703 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_116, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_70, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_139, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_151, S => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_152);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1704 : MAOI222D1BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_145, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_199, C => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_117, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_150);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1705 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_123, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_100, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_126, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_148, S => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_149);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1706 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_67, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_127, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_66, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_146, S => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_147);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1707 : MAOI222D1BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_130, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_135, C => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_110, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_145);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1708 : MAOI222D1BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_131, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_63, C => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_111, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_144);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1709 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_132, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_131, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_132, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_131, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_143);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1710 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_125, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_71, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_120, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_141, S => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_142);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1712 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_128, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_83, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_64, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_138, S => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_139);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1713 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_68, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_91, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_119, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_136, S => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_137);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1714 : MAOI222D1BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_112, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_201, C => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_58, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_135);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1715 : MAOI222D1BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_60, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_114, C => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_77, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_134);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1717 : CKXOR2D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_63, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_111, Z => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_132);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1718 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_115, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_74, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_115, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_74, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_131);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1719 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_59, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_113, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_59, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_113, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_130);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1720 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_122, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_97, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_122, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_97, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_129);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1721 : HA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_102, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_73, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_127, S => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_128);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1722 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_82, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_89, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_86, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_125, S => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_126);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1723 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_84, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_108, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_65, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_123, S => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_124);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1724 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_92, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_93, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_69, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_122, S => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_121);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1725 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_90, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_94, CI => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_85, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_119, S => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_120);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1727 : MAOI222D1BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_59, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_76, C => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_104, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_117);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1728 : MAOI222D1BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_75, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_78, C => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_103, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_116);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1729 : XNR2D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_78, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_103, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_115);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1730 : MOAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_79, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_101, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_79, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_101, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_114);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1731 : CKXOR2D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_76, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_104, Z => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_113);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1732 : MOAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_80, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_107, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_80, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_107, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_112);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1733 : IND2D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_79, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_101, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_111);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1734 : IND2D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_80, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_107, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_110);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1735 : HA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_62, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_72, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_108, S => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_109);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1736 : HA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_95, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_87, CO => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_107, S => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_106);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1737 : OAI21D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_81, A2 => TL02_kb_y_1, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_100, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_105);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1738 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_99, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_93, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_99, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_93, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_104);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1739 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_96, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_98, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_96, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_98, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_103);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1740 : INR2XD0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_98, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_96, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_102);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1741 : INR2D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_99, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_93, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_101);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1742 : ND2D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_81, A2 => TL02_kb_y_1, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_100);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1743 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_94, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_95);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1744 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_91, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_92);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1745 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_89, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_90);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1747 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_55, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_49, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_34, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_99);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1748 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_51, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_33, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_45, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_98);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1749 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_53, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_48, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_36, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_87);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1750 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_23, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_55, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_40, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_34, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_86);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1751 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_40, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_55, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_43, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_34, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_85);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1752 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_47, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_53, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_24, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_36, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_84);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1753 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_20, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_51, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_33, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_97);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1754 : OAI21D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_52, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_32, B => TL02_kb_y_6, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_96);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1755 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_38, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_55, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_42, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_34, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_83);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1756 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_28, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_51, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_15, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_33, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_82);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1757 : OAI21D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_54, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_37, B => TL02_kb_y_3, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_94);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1758 : OAI21D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_56, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_35, B => TL02_kb_y_5, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_93);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1759 : AOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_44, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_56, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_35, B2 => TL02_kb_y_5, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_91);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1760 : AOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_25, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_54, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_37, B2 => TL02_kb_y_3, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_89);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1761 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_74, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_75);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1762 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_18, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_52, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_28, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_33, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_81);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1763 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_51, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_45, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_14, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_33, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_73);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1764 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_16, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_37, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_48, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_53, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_80);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1765 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_22, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_35, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_49, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_55, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_79);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1766 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_14, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_51, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_17, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_33, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_72);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1767 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_15, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_51, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_21, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_33, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_71);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1768 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_41, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_53, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_46, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_36, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_70);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1769 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_19, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_51, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_20, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_33, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_69);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1770 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_22, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_56, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_38, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_34, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_78);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1771 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_27, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_53, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_39, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_36, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_77);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1772 : AOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_16, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_54, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_26, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_37, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_76);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1773 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_21, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_51, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_19, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_33, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_68);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1774 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_42, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_55, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_50, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_34, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_67);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1775 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_46, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_53, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_47, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_36, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_66);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1776 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_39, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_53, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_41, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_36, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_74);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1777 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_50, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_55, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_23, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_34, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_65);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1778 : MOAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_11, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_7, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_8, B2 => TL02_kb_y_0, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_64);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1779 : OA22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_12, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_7, B1 => n_483, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_11, Z => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_63);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1780 : MOAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2, A2 => n_483, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_8, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_6, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_62);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1782 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_10, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_7, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_12, B2 => n_483, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_60);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1783 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_13, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_6, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_10, B2 => n_483, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_59);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1784 : MOAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_9, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_7, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_13, B2 => TL02_kb_y_0, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_58);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1785 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_9, A2 => n_483, B1 => TL02_n_452, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_7, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_57);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1786 : INVD1BWP7T port map(I => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_56, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_55);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1787 : NR2XD0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_31, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_35, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_56);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1788 : INVD1BWP7T port map(I => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_54, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_53);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1789 : NR2XD0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_29, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_37, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_54);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1790 : INVD1BWP7T port map(I => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_52, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_51);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1791 : NR2XD0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_32, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_30, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_52);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1792 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_43, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_44);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1793 : INVD1BWP7T port map(I => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_37, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_36);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1794 : INVD1BWP7T port map(I => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_35, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_34);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1795 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_33, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_32);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1796 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, A2 => TL02_kb_y_4, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, B2 => TL02_kb_y_4, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_31);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1797 : MAOI22D0BWP7T port map(A1 => n_487, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, B1 => n_487, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_30);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1798 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, A2 => TL02_kb_y_2, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, B2 => TL02_kb_y_2, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_29);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1799 : MAOI22D0BWP7T port map(A1 => TL02_n_449, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, B1 => TL02_n_449, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_50);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1800 : MAOI22D0BWP7T port map(A1 => TL02_n_453, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, B1 => TL02_n_453, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_49);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1801 : MAOI22D0BWP7T port map(A1 => TL02_n_453, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, B1 => TL02_n_453, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_48);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1802 : MAOI22D0BWP7T port map(A1 => TL02_n_447, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, B1 => TL02_n_447, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_47);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1803 : MAOI22D0BWP7T port map(A1 => TL02_n_448, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, B1 => TL02_n_448, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_46);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1804 : MAOI22D0BWP7T port map(A1 => TL02_n_453, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, B1 => TL02_n_453, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_45);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1805 : MAOI22D0BWP7T port map(A1 => TL02_n_446, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, B1 => TL02_n_446, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_43);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1806 : MAOI22D0BWP7T port map(A1 => TL02_n_450, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, B1 => TL02_n_450, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_42);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1807 : MAOI22D0BWP7T port map(A1 => TL02_n_449, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, B1 => TL02_n_449, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_41);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1808 : MAOI22D0BWP7T port map(A1 => TL02_n_447, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, B1 => TL02_n_447, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_40);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1809 : MAOI22D0BWP7T port map(A1 => TL02_n_450, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, B1 => TL02_n_450, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_39);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1810 : MAOI22D0BWP7T port map(A1 => TL02_n_451, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, B1 => TL02_n_451, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_38);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1811 : MOAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2, A2 => TL02_kb_y_2, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2, B2 => TL02_kb_y_2, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_37);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1812 : MOAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, A2 => TL02_kb_y_4, B1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, B2 => TL02_kb_y_4, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_35);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1813 : MAOI22D0BWP7T port map(A1 => n_487, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, B1 => n_487, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_33);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1814 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_26, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_27);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1815 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_24, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_25);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1816 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_17, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_18);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1817 : MAOI22D0BWP7T port map(A1 => TL02_n_450, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, B1 => TL02_n_450, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_28);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1818 : MOAI22D0BWP7T port map(A1 => TL02_n_451, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, B1 => TL02_n_451, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_26);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1819 : MAOI22D0BWP7T port map(A1 => TL02_n_446, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, B1 => TL02_n_446, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_24);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1820 : MAOI22D0BWP7T port map(A1 => TL02_n_448, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, B1 => TL02_n_448, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_23);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1821 : MOAI22D0BWP7T port map(A1 => TL02_n_452, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, B1 => TL02_n_452, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_22);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1822 : MAOI22D0BWP7T port map(A1 => TL02_n_448, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, B1 => TL02_n_448, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_21);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1823 : MAOI22D0BWP7T port map(A1 => TL02_n_446, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, B1 => TL02_n_446, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_20);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1824 : MAOI22D0BWP7T port map(A1 => TL02_n_447, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, B1 => TL02_n_447, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_19);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1825 : MAOI22D0BWP7T port map(A1 => TL02_n_451, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, B1 => TL02_n_451, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_17);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1826 : MOAI22D0BWP7T port map(A1 => TL02_n_452, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, B1 => TL02_n_452, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_16);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1827 : MAOI22D0BWP7T port map(A1 => TL02_n_449, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, B1 => TL02_n_449, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_15);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1828 : MAOI22D0BWP7T port map(A1 => TL02_n_452, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, B1 => TL02_n_452, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_14);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1829 : MOAI22D0BWP7T port map(A1 => TL02_n_450, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2, B1 => TL02_n_450, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_13);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1830 : MAOI22D0BWP7T port map(A1 => TL02_n_448, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2, B1 => TL02_n_448, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_12);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1831 : MAOI22D0BWP7T port map(A1 => TL02_n_447, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2, B1 => TL02_n_447, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_11);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1832 : MAOI22D0BWP7T port map(A1 => TL02_n_449, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2, B1 => TL02_n_449, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_10);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1833 : MAOI22D0BWP7T port map(A1 => TL02_n_451, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2, B1 => TL02_n_451, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_9);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1834 : MOAI22D0BWP7T port map(A1 => TL02_n_446, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2, B1 => TL02_n_446, B2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_8);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1835 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_7, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_6);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1836 : CKND2D1BWP7T port map(A1 => n_483, A2 => TL02_kb_y_1, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_7);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1838 : INVD1BWP7T port map(I => TL02_kb_y_6, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_4);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1839 : INVD1BWP7T port map(I => TL02_kb_y_5, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_3);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1840 : INVD1BWP7T port map(I => TL02_kb_y_1, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1841 : INVD1BWP7T port map(I => TL02_kb_y_3, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_1);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g1842 : XOR3D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_114, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_77, A3 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_60, Z => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_199);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g2 : OA21D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_106, A2 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_200, B => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_57, Z => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_201);
  TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_g3 : NR3D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_2, A2 => TL02_n_453, A3 => TL02_n_452, ZN => TL02_PHS1_knockback_mul_36_239_Y_PHS1_knockback_mul_36_97_n_200);
  ATT1_g13365 : NR4D0BWP7T port map(A1 => ATT1_n_759, A2 => ATT1_n_680, A3 => ATT1_n_643, A4 => ATT1_n_638, ZN => dirx1new1(5));
  ATT1_g13366 : NR4D0BWP7T port map(A1 => ATT1_n_758, A2 => ATT1_n_690, A3 => ATT1_n_638, A4 => ATT1_n_630, ZN => dirx1new1(4));
  ATT1_g13367 : IND4D0BWP7T port map(A1 => ATT1_n_690, B1 => ATT1_n_646, B2 => ATT1_n_41, B3 => ATT1_n_757, ZN => ATT1_n_759);
  ATT1_g13368 : MOAI22D0BWP7T port map(A1 => ATT1_n_757, A2 => ATT1_n_738, B1 => ATT1_n_757, B2 => ATT1_n_738, ZN => dirx1new1(6));
  ATT1_g13369 : NR4D0BWP7T port map(A1 => ATT1_n_756, A2 => ATT1_n_681, A3 => ATT1_n_668, A4 => ATT1_n_598, ZN => diry1new1(4));
  ATT1_g13370 : ND4D0BWP7T port map(A1 => ATT1_n_757, A2 => ATT1_n_676, A3 => ATT1_n_42, A4 => ATT1_n_663, ZN => ATT1_n_758);
  ATT1_g13371 : OA21D0BWP7T port map(A1 => ATT1_n_754, A2 => ATT1_n_737, B => ATT1_n_732, Z => diry1new1(7));
  ATT1_g13372 : NR4D0BWP7T port map(A1 => ATT1_n_310, A2 => ATT1_n_755, A3 => ATT1_n_638, A4 => ATT1_n_630, ZN => diry1new1(5));
  ATT1_g13373 : MOAI22D0BWP7T port map(A1 => ATT1_n_753, A2 => ATT1_n_741, B1 => ATT1_n_753, B2 => ATT1_n_741, ZN => dirx1new1(3));
  ATT1_g13374 : CKXOR2D1BWP7T port map(A1 => ATT1_n_754, A2 => ATT1_n_737, Z => diry1new1(6));
  ATT1_g13375 : IND2D1BWP7T port map(A1 => ATT1_n_753, B1 => ATT1_n_741, ZN => ATT1_n_757);
  ATT1_g13376 : ND4D0BWP7T port map(A1 => ATT1_n_754, A2 => ATT1_n_696, A3 => ATT1_n_682, A4 => ATT1_n_652, ZN => ATT1_n_756);
  ATT1_g13377 : ND4D0BWP7T port map(A1 => ATT1_n_754, A2 => ATT1_n_701, A3 => ATT1_n_669, A4 => ATT1_n_586, ZN => ATT1_n_755);
  ATT1_g13378 : MOAI22D0BWP7T port map(A1 => ATT1_n_752, A2 => ATT1_n_743, B1 => ATT1_n_752, B2 => ATT1_n_743, ZN => dirx1new1(2));
  ATT1_g13379 : MOAI22D0BWP7T port map(A1 => ATT1_n_751, A2 => ATT1_n_731, B1 => ATT1_n_751, B2 => ATT1_n_731, ZN => diry1new1(3));
  ATT1_g13380 : IND2D1BWP7T port map(A1 => ATT1_n_751, B1 => ATT1_n_731, ZN => ATT1_n_754);
  ATT1_g13381 : IND2D1BWP7T port map(A1 => ATT1_n_743, B1 => ATT1_n_752, ZN => ATT1_n_753);
  ATT1_g13382 : HA1D0BWP7T port map(A => ATT1_n_712, B => ATT1_n_749, CO => ATT1_n_752, S => dirx1new1(1));
  ATT1_g13383 : MOAI22D0BWP7T port map(A1 => ATT1_n_750, A2 => ATT1_n_739, B1 => ATT1_n_750, B2 => ATT1_n_739, ZN => diry1new1(2));
  ATT1_g13384 : IND2D1BWP7T port map(A1 => ATT1_n_739, B1 => ATT1_n_750, ZN => ATT1_n_751);
  ATT1_g13385 : HA1D0BWP7T port map(A => ATT1_n_735, B => ATT1_n_746, CO => ATT1_n_750, S => diry1new1(1));
  ATT1_g13386 : ND4D0BWP7T port map(A1 => ATT1_n_747, A2 => ATT1_n_636, A3 => ATT1_n_625, A4 => ATT1_n_472, ZN => dirx2new1(0));
  ATT1_g13387 : INVD1BWP7T port map(I => dirx1new1(0), ZN => ATT1_n_749);
  ATT1_g13388 : OAI211D1BWP7T port map(A1 => ATT1_n_489, A2 => ATT1_n_431, B => ATT1_n_748, C => ATT1_n_458, ZN => dirx1new1(0));
  ATT1_g13389 : AOI222D0BWP7T port map(A1 => ATT1_n_745, A2 => ATT1_n_697, B1 => ATT1_n_530, B2 => ATT1_n_540, C1 => ATT1_n_512, C2 => ATT1_n_592, ZN => ATT1_n_748);
  ATT1_g13390 : OA32D1BWP7T port map(A1 => ATT1_n_479, A2 => ATT1_n_744, A3 => FE_OFN2_ATT1_n_301, B1 => ATT1_n_493, B2 => ATT1_n_431, Z => ATT1_n_747);
  ATT1_g13391 : INVD0BWP7T port map(I => ATT1_n_746, ZN => diry1new1(0));
  ATT1_g13392 : AOI221D1BWP7T port map(A1 => ATT1_n_361, A2 => ATT1_n_742, B1 => ATT1_n_512, B2 => ATT1_n_451, C => ATT1_n_664, ZN => ATT1_n_746);
  ATT1_g13393 : NR4D0BWP7T port map(A1 => ATT1_n_740, A2 => ATT1_n_605, A3 => ATT1_n_601, A4 => ATT1_n_513, ZN => ATT1_n_745);
  ATT1_g13394 : ND4D0BWP7T port map(A1 => ATT1_n_316, A2 => ATT1_n_736, A3 => ATT1_n_523, A4 => ATT1_n_493, ZN => ATT1_n_744);
  ATT1_g13395 : OR4D1BWP7T port map(A1 => ATT1_n_630, A2 => ATT1_n_643, A3 => ATT1_n_667, A4 => ATT1_n_730, Z => ATT1_n_743);
  ATT1_g13396 : NR4D0BWP7T port map(A1 => ATT1_n_733, A2 => ATT1_n_648, A3 => ATT1_n_680, A4 => ATT1_n_667, ZN => ATT1_n_742);
  ATT1_g13397 : NR4D0BWP7T port map(A1 => ATT1_n_728, A2 => ATT1_n_681, A3 => ATT1_n_680, A4 => ATT1_n_668, ZN => ATT1_n_741);
  ATT1_g13398 : OAI211D1BWP7T port map(A1 => ATT1_n_521, A2 => ATT1_n_364, B => ATT1_n_734, C => ATT1_n_682, ZN => ATT1_n_740);
  ATT1_g13399 : ND4D0BWP7T port map(A1 => ATT1_n_724, A2 => ATT1_n_642, A3 => ATT1_n_647, A4 => ATT1_n_641, ZN => dirx2new1(4));
  ATT1_g13400 : ND3D0BWP7T port map(A1 => ATT1_n_727, A2 => ATT1_n_480, A3 => ATT1_n_490, ZN => dirx2new1(6));
  ATT1_g13401 : ND4D0BWP7T port map(A1 => ATT1_n_725, A2 => ATT1_n_640, A3 => ATT1_n_641, A4 => ATT1_n_599, ZN => dirx2new1(2));
  ATT1_g13402 : ND4D0BWP7T port map(A1 => ATT1_n_723, A2 => ATT1_n_640, A3 => ATT1_n_641, A4 => ATT1_n_550, ZN => diry2new1(4));
  ATT1_g13403 : ND4D0BWP7T port map(A1 => ATT1_n_726, A2 => ATT1_n_647, A3 => ATT1_n_597, A4 => ATT1_n_550, ZN => diry2new1(3));
  ATT1_g13404 : IND4D0BWP7T port map(A1 => ATT1_n_680, B1 => ATT1_n_639, B2 => ATT1_n_697, B3 => ATT1_n_719, ZN => ATT1_n_739);
  ATT1_g13405 : ND4D0BWP7T port map(A1 => ATT1_n_721, A2 => ATT1_n_645, A3 => ATT1_n_644, A4 => ATT1_n_651, ZN => diry2new1(0));
  ATT1_g13406 : ND4D0BWP7T port map(A1 => ATT1_n_720, A2 => ATT1_n_670, A3 => ATT1_n_641, A4 => ATT1_n_597, ZN => diry2new1(2));
  ATT1_g13407 : AN4D0BWP7T port map(A1 => ATT1_n_718, A2 => ATT1_n_558, A3 => ATT1_n_526, A4 => ATT1_n_817, Z => ATT1_n_736);
  ATT1_g13408 : NR4D0BWP7T port map(A1 => ATT1_n_717, A2 => ATT1_n_499, A3 => ATT1_n_451, A4 => ATT1_n_467, ZN => ATT1_n_738);
  ATT1_g13409 : OAI21D0BWP7T port map(A1 => ATT1_n_456, A2 => ATT1_n_559, B => ATT1_n_732, ZN => ATT1_n_737);
  ATT1_g13410 : AN3D1BWP7T port map(A1 => ATT1_n_729, A2 => ATT1_n_697, A3 => ATT1_n_639, Z => ATT1_n_735);
  ATT1_g13411 : INVD0BWP7T port map(I => ATT1_n_733, ZN => ATT1_n_734);
  ATT1_g13412 : ND4D0BWP7T port map(A1 => ATT1_n_715, A2 => ATT1_n_642, A3 => ATT1_n_640, A4 => ATT1_n_644, ZN => dirx2new1(5));
  ATT1_g13413 : ND3D0BWP7T port map(A1 => ATT1_n_722, A2 => ATT1_n_559, A3 => ATT1_n_496, ZN => ATT1_n_733);
  ATT1_g13414 : IND4D0BWP7T port map(A1 => ATT1_n_385, B1 => ATT1_n_697, B2 => ATT1_n_709, B3 => ATT1_n_320, ZN => ATT1_n_732);
  ATT1_g13415 : NR4D0BWP7T port map(A1 => ATT1_n_710, A2 => ATT1_n_681, A3 => ATT1_n_680, A4 => ATT1_n_601, ZN => ATT1_n_731);
  ATT1_g13416 : IND4D0BWP7T port map(A1 => ATT1_n_648, B1 => ATT1_n_612, B2 => ATT1_n_646, B3 => ATT1_n_716, ZN => ATT1_n_730);
  ATT1_g13417 : ND4D0BWP7T port map(A1 => ATT1_n_714, A2 => ATT1_n_698, A3 => ATT1_n_649, A4 => ATT1_n_644, ZN => diry2new1(1));
  ATT1_g13418 : ND4D0BWP7T port map(A1 => ATT1_n_711, A2 => ATT1_n_698, A3 => ATT1_n_642, A4 => ATT1_n_599, ZN => dirx2new1(3));
  ATT1_g13419 : ND4D0BWP7T port map(A1 => ATT1_n_713, A2 => ATT1_n_642, A3 => ATT1_n_640, A4 => ATT1_n_600, ZN => diry2new1(5));
  ATT1_g13420 : NR4D0BWP7T port map(A1 => ATT1_n_703, A2 => ATT1_n_668, A3 => ATT1_n_601, A4 => ATT1_n_513, ZN => ATT1_n_729);
  ATT1_g13421 : OR4D1BWP7T port map(A1 => ATT1_n_513, A2 => ATT1_n_643, A3 => ATT1_n_690, A4 => ATT1_n_704, Z => ATT1_n_728);
  ATT1_g13422 : AN4D0BWP7T port map(A1 => ATT1_n_699, A2 => ATT1_n_649, A3 => ATT1_n_600, A4 => ATT1_n_533, Z => ATT1_n_727);
  ATT1_g13423 : AN3D0BWP7T port map(A1 => ATT1_n_700, A2 => ATT1_n_670, A3 => ATT1_n_651, Z => ATT1_n_726);
  ATT1_g13424 : AN4D0BWP7T port map(A1 => ATT1_n_695, A2 => ATT1_n_645, A3 => ATT1_n_644, A4 => ATT1_n_597, Z => ATT1_n_725);
  ATT1_g13425 : NR2XD0BWP7T port map(A1 => ATT1_n_691, A2 => ATT1_n_708, ZN => ATT1_n_724);
  ATT1_g13426 : AN3D0BWP7T port map(A1 => ATT1_n_702, A2 => ATT1_n_651, A3 => ATT1_n_602, Z => ATT1_n_723);
  ATT1_g13427 : NR3D0BWP7T port map(A1 => ATT1_n_385, A2 => ATT1_n_706, A3 => ATT1_n_534, ZN => ATT1_n_722);
  ATT1_g13428 : NR4D0BWP7T port map(A1 => ATT1_n_689, A2 => ATT1_n_693, A3 => ATT1_n_650, A4 => ATT1_n_607, ZN => ATT1_n_721);
  ATT1_g13429 : NR4D0BWP7T port map(A1 => ATT1_n_683, A2 => ATT1_n_689, A3 => ATT1_n_694, A4 => ATT1_n_603, ZN => ATT1_n_720);
  ATT1_g13430 : NR2XD0BWP7T port map(A1 => ATT1_n_707, A2 => ATT1_n_667, ZN => ATT1_n_719);
  ATT1_g13431 : AN4D0BWP7T port map(A1 => ATT1_n_688, A2 => ATT1_n_661, A3 => ATT1_n_599, A4 => ATT1_n_600, Z => ATT1_n_718);
  ATT1_g13432 : ND4D0BWP7T port map(A1 => ATT1_n_686, A2 => ATT1_n_632, A3 => ATT1_n_604, A4 => ATT1_n_539, ZN => ATT1_n_717);
  ATT1_g13433 : AN4D0BWP7T port map(A1 => ATT1_n_677, A2 => ATT1_n_631, A3 => ATT1_n_637, A4 => ATT1_n_458, Z => ATT1_n_716);
  ATT1_g13434 : AN4D0BWP7T port map(A1 => ATT1_n_698, A2 => ATT1_n_692, A3 => ATT1_n_684, A4 => ATT1_n_675, Z => ATT1_n_715);
  ATT1_g13436 : NR4D0BWP7T port map(A1 => ATT1_n_683, A2 => ATT1_n_665, A3 => ATT1_n_666, A4 => ATT1_n_487, ZN => ATT1_n_714);
  ATT1_g13437 : INR4D0BWP7T port map(A1 => ATT1_n_670, B1 => ATT1_n_655, B2 => ATT1_n_674, B3 => ATT1_n_683, ZN => ATT1_n_713);
  ATT1_g13438 : NR4D0BWP7T port map(A1 => ATT1_n_648, A2 => ATT1_n_679, A3 => ATT1_n_638, A4 => ATT1_n_598, ZN => ATT1_n_712);
  ATT1_g13439 : AN4D0BWP7T port map(A1 => ATT1_n_692, A2 => ATT1_n_678, A3 => ATT1_n_635, A4 => ATT1_n_602, Z => ATT1_n_711);
  ATT1_g13440 : IND4D0BWP7T port map(A1 => ATT1_n_598, B1 => ATT1_n_604, B2 => ATT1_n_669, B3 => ATT1_n_673, ZN => ATT1_n_710);
  ATT1_g13441 : OAI21D0BWP7T port map(A1 => ATT1_n_671, A2 => ATT1_n_412, B => ATT1_n_706, ZN => ATT1_n_709);
  ATT1_g13442 : IND4D0BWP7T port map(A1 => ATT1_n_691, B1 => ATT1_n_599, B2 => ATT1_n_628, B3 => ATT1_n_584, ZN => dirx2new1(1));
  ATT1_g13443 : OAI211D1BWP7T port map(A1 => ATT1_n_480, A2 => ATT1_n_483, B => ATT1_n_687, C => ATT1_n_575, ZN => ATT1_n_708);
  ATT1_g13444 : ND4D0BWP7T port map(A1 => ATT1_n_658, A2 => ATT1_n_669, A3 => ATT1_n_646, A4 => ATT1_n_569, ZN => ATT1_n_707);
  ATT1_g13445 : IND4D0BWP7T port map(A1 => ATT1_n_668, B1 => ATT1_n_633, B2 => ATT1_n_42, B3 => ATT1_n_634, ZN => ATT1_n_705);
  ATT1_g13446 : OAI211D1BWP7T port map(A1 => ATT1_n_508, A2 => ATT1_n_447, B => ATT1_n_672, C => ATT1_n_543, ZN => ATT1_n_704);
  ATT1_g13447 : ND4D0BWP7T port map(A1 => ATT1_n_589, A2 => ATT1_n_613, A3 => ATT1_n_660, A4 => ATT1_n_611, ZN => ATT1_n_703);
  ATT1_g13448 : IND3D1BWP7T port map(A1 => ATT1_n_671, B1 => ATT1_n_316, B2 => ATT1_n_347, ZN => ATT1_n_706);
  ATT1_g13449 : NR4D0BWP7T port map(A1 => ATT1_n_685, A2 => ATT1_n_616, A3 => ATT1_n_629, A4 => ATT1_n_564, ZN => ATT1_n_702);
  ATT1_g13450 : INR3D0BWP7T port map(A1 => ATT1_n_682, B1 => ATT1_n_605, B2 => ATT1_n_626, ZN => ATT1_n_701);
  ATT1_g13451 : NR4D0BWP7T port map(A1 => ATT1_n_617, A2 => ATT1_n_603, A3 => ATT1_n_606, A4 => ATT1_n_570, ZN => ATT1_n_700);
  ATT1_g13452 : AOI22D0BWP7T port map(A1 => FE_OFN2_ATT1_n_301, A2 => ATT1_n_662, B1 => ATT1_n_352, B2 => ATT1_n_470, ZN => ATT1_n_699);
  ATT1_g13453 : NR3D0BWP7T port map(A1 => ATT1_n_657, A2 => ATT1_n_580, A3 => ATT1_n_546, ZN => ATT1_n_696);
  ATT1_g13454 : NR4D0BWP7T port map(A1 => ATT1_n_623, A2 => ATT1_n_591, A3 => ATT1_n_572, A4 => ATT1_n_590, ZN => ATT1_n_695);
  ATT1_g13455 : OAI221D0BWP7T port map(A1 => ATT1_n_517, A2 => ATT1_n_531, B1 => ATT1_n_480, B2 => ATT1_n_407, C => ATT1_n_656, ZN => ATT1_n_694);
  ATT1_g13456 : OAI221D0BWP7T port map(A1 => ATT1_n_443, A2 => ATT1_n_558, B1 => ATT1_n_526, B2 => ATT1_n_434, C => ATT1_n_659, ZN => ATT1_n_693);
  ATT1_g13457 : NR2XD0BWP7T port map(A1 => ATT1_n_685, A2 => ATT1_n_603, ZN => ATT1_n_698);
  ATT1_g13458 : NR2D1BWP7T port map(A1 => ATT1_n_681, A2 => ATT1_n_653, ZN => ATT1_n_697);
  ATT1_g13459 : CKND1BWP7T port map(I => ATT1_n_689, ZN => ATT1_n_688);
  ATT1_g13460 : NR4D0BWP7T port map(A1 => ATT1_n_620, A2 => ATT1_n_552, A3 => ATT1_n_545, A4 => ATT1_n_588, ZN => ATT1_n_687);
  ATT1_g13461 : AOI211XD0BWP7T port map(A1 => ATT1_n_317, A2 => ATT1_n_412, B => ATT1_n_624, C => ATT1_n_653, ZN => ATT1_n_686);
  ATT1_g13462 : OA211D0BWP7T port map(A1 => ATT1_n_560, A2 => ATT1_n_400, B => ATT1_n_641, C => ATT1_n_645, Z => ATT1_n_692);
  ATT1_g13463 : OAI21D0BWP7T port map(A1 => ATT1_n_422, A2 => ATT1_n_441, B => ATT1_n_684, ZN => ATT1_n_691);
  ATT1_g13464 : AO211D0BWP7T port map(A1 => ATT1_n_399, A2 => ATT1_n_439, B => ATT1_n_667, C => ATT1_n_605, Z => ATT1_n_690);
  ATT1_g13465 : ND3D0BWP7T port map(A1 => ATT1_n_647, A2 => ATT1_n_649, A3 => ATT1_n_640, ZN => ATT1_n_689);
  ATT1_g13466 : ND3D0BWP7T port map(A1 => ATT1_n_565, A2 => ATT1_n_563, A3 => ATT1_n_579, ZN => ATT1_n_679);
  ATT1_g13467 : OA221D0BWP7T port map(A1 => ATT1_n_390, A2 => ATT1_n_560, B1 => ATT1_n_438, B2 => ATT1_n_477, C => ATT1_n_582, Z => ATT1_n_678);
  ATT1_g13468 : AOI221D0BWP7T port map(A1 => ATT1_n_453, A2 => ATT1_n_488, B1 => ATT1_n_532, B2 => ATT1_n_451, C => ATT1_n_618, ZN => ATT1_n_677);
  ATT1_g13469 : AOI211XD0BWP7T port map(A1 => ATT1_n_378, A2 => ATT1_n_39, B => ATT1_n_567, C => ATT1_n_583, ZN => ATT1_n_676);
  ATT1_g13470 : NR4D0BWP7T port map(A1 => ATT1_n_585, A2 => ATT1_n_578, A3 => ATT1_n_576, A4 => ATT1_n_505, ZN => ATT1_n_675);
  ATT1_g13471 : OAI221D0BWP7T port map(A1 => ATT1_n_433, A2 => ATT1_n_561, B1 => ATT1_n_480, B2 => ATT1_n_455, C => ATT1_n_619, ZN => ATT1_n_674);
  ATT1_g13472 : AOI221D0BWP7T port map(A1 => ATT1_n_519, A2 => ATT1_n_482, B1 => ATT1_n_387, B2 => ATT1_n_451, C => ATT1_n_621, ZN => ATT1_n_673);
  ATT1_g13473 : OA221D0BWP7T port map(A1 => ATT1_n_415, A2 => ATT1_n_539, B1 => ATT1_n_442, B2 => ATT1_n_445, C => ATT1_n_627, Z => ATT1_n_672);
  ATT1_g13474 : IND2D1BWP7T port map(A1 => ATT1_n_655, B1 => ATT1_n_647, ZN => ATT1_n_685);
  ATT1_g13476 : NR2XD0BWP7T port map(A1 => ATT1_n_650, A2 => ATT1_n_610, ZN => ATT1_n_684);
  ATT1_g13477 : IND2D1BWP7T port map(A1 => ATT1_n_650, B1 => ATT1_n_550, ZN => ATT1_n_683);
  ATT1_g13478 : AN2D1BWP7T port map(A1 => ATT1_n_646, A2 => ATT1_n_604, Z => ATT1_n_682);
  ATT1_g13479 : CKND2D1BWP7T port map(A1 => ATT1_n_586, A2 => ATT1_n_654, ZN => ATT1_n_681);
  ATT1_g13480 : IND2D1BWP7T port map(A1 => ATT1_n_630, B1 => ATT1_n_611, ZN => ATT1_n_680);
  ATT1_g13481 : OAI22D0BWP7T port map(A1 => ATT1_n_609, A2 => ATT1_n_480, B1 => ATT1_n_38, B2 => ATT1_n_523, ZN => ATT1_n_666);
  ATT1_g13482 : OAI221D0BWP7T port map(A1 => ATT1_n_426, A2 => ATT1_n_561, B1 => ATT1_n_526, B2 => ATT1_n_367, C => ATT1_n_615, ZN => ATT1_n_665);
  ATT1_g13483 : OAI221D0BWP7T port map(A1 => ATT1_n_460, A2 => ATT1_n_496, B1 => ATT1_n_489, B2 => ATT1_n_461, C => ATT1_n_622, ZN => ATT1_n_664);
  ATT1_g13484 : AOI221D0BWP7T port map(A1 => ATT1_n_562, A2 => ATT1_n_488, B1 => ATT1_n_529, B2 => ATT1_n_439, C => ATT1_n_506, ZN => ATT1_n_663);
  ATT1_g13485 : ND4D0BWP7T port map(A1 => ATT1_n_555, A2 => ATT1_n_560, A3 => ATT1_n_510, A4 => ATT1_n_441, ZN => ATT1_n_662);
  ATT1_g13486 : AOI211XD0BWP7T port map(A1 => ATT1_n_360, A2 => ATT1_n_528, B => ATT1_n_606, C => ATT1_n_607, ZN => ATT1_n_661);
  ATT1_g13487 : AOI22D0BWP7T port map(A1 => ATT1_n_608, A2 => ATT1_n_451, B1 => ATT1_n_366, B2 => ATT1_n_482, ZN => ATT1_n_660);
  ATT1_g13488 : AOI21D0BWP7T port map(A1 => ATT1_n_512, A2 => ATT1_n_479, B => ATT1_n_614, ZN => ATT1_n_659);
  ATT1_g13489 : AOI31D0BWP7T port map(A1 => ATT1_n_551, A2 => ATT1_n_309, A3 => ATT1_n_497, B => ATT1_n_573, ZN => ATT1_n_658);
  ATT1_g13490 : OAI222D0BWP7T port map(A1 => ATT1_n_409, A2 => ATT1_n_559, B1 => ATT1_n_489, B2 => ATT1_n_410, C1 => ATT1_n_521, C2 => ATT1_n_435, ZN => ATT1_n_657);
  ATT1_g13491 : AOI31D0BWP7T port map(A1 => ATT1_n_551, A2 => ATT1_n_309, A3 => ATT1_n_524, B => ATT1_n_587, ZN => ATT1_n_656);
  ATT1_g13492 : IOA21D1BWP7T port map(A1 => ATT1_n_358, A2 => orientationp2, B => ATT1_n_632, ZN => ATT1_n_671);
  ATT1_g13493 : OA21D0BWP7T port map(A1 => ATT1_n_416, A2 => ATT1_n_558, B => ATT1_n_645, Z => ATT1_n_670);
  ATT1_g13494 : IAO21D0BWP7T port map(A1 => ATT1_n_416, A2 => ATT1_n_559, B => ATT1_n_643, ZN => ATT1_n_669);
  ATT1_g13495 : IOA21D1BWP7T port map(A1 => ATT1_n_310, A2 => ATT1_n_596, B => ATT1_n_612, ZN => ATT1_n_668);
  ATT1_g13496 : OAI21D0BWP7T port map(A1 => ATT1_n_376, A2 => ATT1_n_521, B => ATT1_n_652, ZN => ATT1_n_667);
  ATT1_g13498 : INVD1BWP7T port map(I => ATT1_n_639, ZN => ATT1_n_638);
  ATT1_g13499 : AOI221D0BWP7T port map(A1 => ATT1_n_512, A2 => ATT1_n_439, B1 => ATT1_n_394, B2 => ATT1_n_467, C => ATT1_n_574, ZN => ATT1_n_637);
  ATT1_g13500 : CKND2D1BWP7T port map(A1 => ATT1_n_530, A2 => ATT1_n_566, ZN => ATT1_n_636);
  ATT1_g13501 : OA221D0BWP7T port map(A1 => ATT1_n_415, A2 => ATT1_n_533, B1 => ATT1_n_510, B2 => ATT1_n_447, C => ATT1_n_581, Z => ATT1_n_635);
  ATT1_g13502 : AOI221D0BWP7T port map(A1 => ATT1_n_383, A2 => ATT1_n_522, B1 => ATT1_n_405, B2 => ATT1_n_499, C => ATT1_n_504, ZN => ATT1_n_634);
  ATT1_g13503 : AOI221D0BWP7T port map(A1 => ATT1_n_514, A2 => ATT1_n_488, B1 => ATT1_n_382, B2 => ATT1_n_39, C => ATT1_n_542, ZN => ATT1_n_633);
  ATT1_g13504 : AN2D1BWP7T port map(A1 => ATT1_n_310, A2 => ATT1_n_595, Z => ATT1_n_655);
  ATT1_g13505 : ND2D1BWP7T port map(A1 => ATT1_n_373, A2 => ATT1_n_596, ZN => ATT1_n_654);
  ATT1_g13506 : INR2XD0BWP7T port map(A1 => ATT1_n_596, B1 => ATT1_n_376, ZN => ATT1_n_653);
  ATT1_g13507 : ND2D1BWP7T port map(A1 => ATT1_n_368, A2 => ATT1_n_596, ZN => ATT1_n_652);
  ATT1_g13508 : INR2XD0BWP7T port map(A1 => ATT1_n_600, B1 => ATT1_n_610, ZN => ATT1_n_651);
  ATT1_g13509 : NR2D1BWP7T port map(A1 => ATT1_n_375, A2 => ATT1_n_594, ZN => ATT1_n_650);
  ATT1_g13510 : IND2D1BWP7T port map(A1 => ATT1_n_376, B1 => ATT1_n_595, ZN => ATT1_n_649);
  ATT1_g13511 : IND2D1BWP7T port map(A1 => ATT1_n_513, B1 => ATT1_n_586, ZN => ATT1_n_648);
  ATT1_g13512 : CKND2D1BWP7T port map(A1 => ATT1_n_373, A2 => ATT1_n_595, ZN => ATT1_n_647);
  ATT1_g13513 : ND2D1BWP7T port map(A1 => ATT1_n_424, A2 => ATT1_n_596, ZN => ATT1_n_646);
  ATT1_g13514 : IND2D1BWP7T port map(A1 => ATT1_n_309, B1 => ATT1_n_595, ZN => ATT1_n_645);
  ATT1_g13515 : INR2XD0BWP7T port map(A1 => ATT1_n_602, B1 => ATT1_n_606, ZN => ATT1_n_644);
  ATT1_g13516 : INR2D1BWP7T port map(A1 => ATT1_n_596, B1 => ATT1_n_309, ZN => ATT1_n_643);
  ATT1_g13517 : INR2XD0BWP7T port map(A1 => ATT1_n_597, B1 => ATT1_n_607, ZN => ATT1_n_642);
  ATT1_g13518 : CKND2D1BWP7T port map(A1 => ATT1_n_368, A2 => ATT1_n_595, ZN => ATT1_n_641);
  ATT1_g13519 : CKND2D1BWP7T port map(A1 => ATT1_n_424, A2 => ATT1_n_595, ZN => ATT1_n_640);
  ATT1_g13520 : CKND2D1BWP7T port map(A1 => ATT1_n_374, A2 => ATT1_n_596, ZN => ATT1_n_639);
  ATT1_g13522 : OAI22D0BWP7T port map(A1 => ATT1_n_409, A2 => ATT1_n_558, B1 => ATT1_n_516, B2 => ATT1_n_480, ZN => ATT1_n_629);
  ATT1_g13523 : AOI221D0BWP7T port map(A1 => ATT1_n_532, A2 => ATT1_n_501, B1 => ATT1_n_403, B2 => ATT1_n_491, C => ATT1_n_568, ZN => ATT1_n_628);
  ATT1_g13524 : AOI211XD0BWP7T port map(A1 => ATT1_n_462, A2 => ATT1_n_451, B => ATT1_n_571, C => ATT1_n_554, ZN => ATT1_n_627);
  ATT1_g13525 : OAI21D0BWP7T port map(A1 => ATT1_n_456, A2 => ATT1_n_558, B => ATT1_n_518, ZN => diry2new1(6));
  ATT1_g13526 : OAI211D1BWP7T port map(A1 => ATT1_n_450, A2 => ATT1_n_455, B => ATT1_n_577, C => ATT1_n_547, ZN => ATT1_n_626);
  ATT1_g13527 : NR3D0BWP7T port map(A1 => ATT1_n_553, A2 => ATT1_n_451, A3 => ATT1_n_467, ZN => dirx1new1(7));
  ATT1_g13528 : IOA21D0BWP7T port map(A1 => ATT1_n_558, A2 => ATT1_n_490, B => ATT1_n_512, ZN => ATT1_n_625);
  ATT1_g13529 : AOI31D0BWP7T port map(A1 => ATT1_n_521, A2 => ATT1_n_508, A3 => ATT1_n_471, B => ATT1_n_300, ZN => ATT1_n_624);
  ATT1_g13530 : OAI211D1BWP7T port map(A1 => ATT1_n_438, A2 => ATT1_n_511, B => ATT1_n_541, C => ATT1_n_472, ZN => ATT1_n_623);
  ATT1_g13531 : ND4D0BWP7T port map(A1 => ATT1_n_533, A2 => ATT1_n_480, A3 => ATT1_n_495, A4 => ATT1_n_490, ZN => dirx2new1(7));
  ATT1_g13532 : OA22D0BWP7T port map(A1 => ATT1_n_443, A2 => ATT1_n_559, B1 => ATT1_n_481, B2 => ATT1_n_434, Z => ATT1_n_622);
  ATT1_g13533 : OAI222D0BWP7T port map(A1 => ATT1_n_437, A2 => ATT1_n_521, B1 => ATT1_n_496, B2 => ATT1_n_537, C1 => ATT1_n_489, C2 => ATT1_n_459, ZN => ATT1_n_621);
  ATT1_g13534 : OAI31D0BWP7T port map(A1 => ATT1_n_495, A2 => FE_OFN2_ATT1_n_301, A3 => ATT1_n_378, B => ATT1_n_593, ZN => ATT1_n_620);
  ATT1_g13535 : OA222D0BWP7T port map(A1 => ATT1_n_452, A2 => ATT1_n_531, B1 => ATT1_n_523, B2 => ATT1_n_408, C1 => ATT1_n_526, C2 => ATT1_n_486, Z => ATT1_n_619);
  ATT1_g13536 : OAI32D1BWP7T port map(A1 => ATT1_n_508, A2 => FE_OFN2_ATT1_n_301, A3 => ATT1_n_391, B1 => ATT1_n_498, B2 => ATT1_n_414, ZN => ATT1_n_618);
  ATT1_g13537 : OAI221D0BWP7T port map(A1 => ATT1_n_537, A2 => ATT1_n_523, B1 => ATT1_n_531, B2 => ATT1_n_459, C => ATT1_n_503, ZN => ATT1_n_617);
  ATT1_g13538 : OAI222D0BWP7T port map(A1 => ATT1_n_410, A2 => ATT1_n_531, B1 => ATT1_n_40, B2 => ATT1_n_435, C1 => ATT1_n_526, C2 => ATT1_n_455, ZN => ATT1_n_616);
  ATT1_g13539 : OA22D0BWP7T port map(A1 => ATT1_n_477, A2 => ATT1_n_531, B1 => ATT1_n_558, B2 => ATT1_n_420, Z => ATT1_n_615);
  ATT1_g13540 : OAI22D0BWP7T port map(A1 => ATT1_n_461, A2 => ATT1_n_561, B1 => ATT1_n_460, B2 => ATT1_n_523, ZN => ATT1_n_614);
  ATT1_g13541 : OA22D0BWP7T port map(A1 => ATT1_n_420, A2 => ATT1_n_559, B1 => ATT1_n_496, B2 => ATT1_n_38, Z => ATT1_n_613);
  ATT1_g13542 : AOI22D0BWP7T port map(A1 => FE_OFN2_ATT1_n_301, A2 => ATT1_n_556, B1 => ATT1_n_317, B2 => ATT1_n_425, ZN => ATT1_n_632);
  ATT1_g13543 : AOI21D0BWP7T port map(A1 => ATT1_n_378, A2 => ATT1_n_522, B => ATT1_n_601, ZN => ATT1_n_631);
  ATT1_g13544 : OAI222D0BWP7T port map(A1 => ATT1_n_349, A2 => ATT1_n_557, B1 => ATT1_n_502, B2 => ATT1_n_332, C1 => ATT1_n_444, C2 => ATT1_n_353, ZN => ATT1_n_630);
  ATT1_g13545 : INVD0BWP7T port map(I => ATT1_n_608, ZN => ATT1_n_609);
  ATT1_g13546 : INVD0BWP7T port map(I => ATT1_n_595, ZN => ATT1_n_594);
  ATT1_g13547 : IND2D1BWP7T port map(A1 => ATT1_n_493, B1 => ATT1_n_562, ZN => ATT1_n_593);
  ATT1_g13548 : ND2D1BWP7T port map(A1 => ATT1_n_559, A2 => ATT1_n_466, ZN => ATT1_n_592);
  ATT1_g13549 : OAI21D0BWP7T port map(A1 => ATT1_n_414, A2 => ATT1_n_495, B => ATT1_n_544, ZN => ATT1_n_591);
  ATT1_g13550 : NR3D0BWP7T port map(A1 => ATT1_n_391, A2 => FE_OFN2_ATT1_n_301, A3 => ATT1_n_510, ZN => ATT1_n_590);
  ATT1_g13551 : MAOI22D0BWP7T port map(A1 => ATT1_n_520, A2 => ATT1_n_488, B1 => ATT1_n_426, B2 => ATT1_n_521, ZN => ATT1_n_589);
  ATT1_g13552 : AOI21D0BWP7T port map(A1 => ATT1_n_530, A2 => ATT1_n_400, B => ATT1_n_438, ZN => ATT1_n_588);
  ATT1_g13553 : OAI22D0BWP7T port map(A1 => ATT1_n_538, A2 => ATT1_n_526, B1 => ATT1_n_436, B2 => ATT1_n_40, ZN => ATT1_n_587);
  ATT1_g13554 : CKND2D1BWP7T port map(A1 => ATT1_n_343, A2 => ATT1_n_556, ZN => ATT1_n_612);
  ATT1_g13555 : ND2D1BWP7T port map(A1 => ATT1_n_337, A2 => ATT1_n_556, ZN => ATT1_n_611);
  ATT1_g13556 : NR2D1BWP7T port map(A1 => ATT1_n_318, A2 => ATT1_n_555, ZN => ATT1_n_610);
  ATT1_g13557 : NR3D0BWP7T port map(A1 => ATT1_n_507, A2 => ATT1_n_368, A3 => FE_OFN2_ATT1_n_301, ZN => ATT1_n_608);
  ATT1_g13558 : NR2D1BWP7T port map(A1 => ATT1_n_324, A2 => ATT1_n_555, ZN => ATT1_n_607);
  ATT1_g13559 : NR2D1BWP7T port map(A1 => ATT1_n_336, A2 => ATT1_n_555, ZN => ATT1_n_606);
  ATT1_g13560 : NR2XD0BWP7T port map(A1 => ATT1_n_324, A2 => ATT1_n_557, ZN => ATT1_n_605);
  ATT1_g13561 : ND2D1BWP7T port map(A1 => ATT1_n_331, A2 => ATT1_n_556, ZN => ATT1_n_604);
  ATT1_g13562 : NR2D1BWP7T port map(A1 => ATT1_n_338, A2 => ATT1_n_555, ZN => ATT1_n_603);
  ATT1_g13563 : IND2D1BWP7T port map(A1 => ATT1_n_555, B1 => ATT1_n_343, ZN => ATT1_n_602);
  ATT1_g13564 : NR2XD0BWP7T port map(A1 => ATT1_n_336, A2 => ATT1_n_557, ZN => ATT1_n_601);
  ATT1_g13565 : OR2D1BWP7T port map(A1 => ATT1_n_332, A2 => ATT1_n_555, Z => ATT1_n_600);
  ATT1_g13566 : AOI211XD0BWP7T port map(A1 => ATT1_n_478, A2 => ATT1_n_430, B => ATT1_n_549, C => ATT1_n_487, ZN => ATT1_n_599);
  ATT1_g13567 : NR2D1BWP7T port map(A1 => ATT1_n_318, A2 => ATT1_n_557, ZN => ATT1_n_598);
  ATT1_g13568 : OR2D1BWP7T port map(A1 => ATT1_n_349, A2 => ATT1_n_555, Z => ATT1_n_597);
  ATT1_g13569 : NR2XD0BWP7T port map(A1 => ATT1_n_417, A2 => ATT1_n_557, ZN => ATT1_n_596);
  ATT1_g13570 : NR2D1BWP7T port map(A1 => ATT1_n_417, A2 => ATT1_n_555, ZN => ATT1_n_595);
  ATT1_g13571 : AO22D0BWP7T port map(A1 => ATT1_n_383, A2 => ATT1_n_528, B1 => ATT1_n_494, B2 => ATT1_n_405, Z => ATT1_n_585);
  ATT1_g13572 : AOI222D0BWP7T port map(A1 => ATT1_n_364, A2 => ATT1_n_492, B1 => ATT1_n_397, B2 => ATT1_n_479, C1 => ATT1_n_355, C2 => ATT1_n_509, ZN => ATT1_n_584);
  ATT1_g13573 : OAI32D0BWP7T port map(A1 => ATT1_n_468, A2 => ATT1_n_484, A3 => ATT1_n_478, B1 => ATT1_n_450, B2 => ATT1_n_483, ZN => ATT1_n_583);
  ATT1_g13574 : AOI21D0BWP7T port map(A1 => ATT1_n_462, A2 => ATT1_n_479, B => ATT1_n_548, ZN => ATT1_n_582);
  ATT1_g13575 : MAOI22D0BWP7T port map(A1 => ATT1_n_535, A2 => ATT1_n_491, B1 => ATT1_n_445, B2 => ATT1_n_441, ZN => ATT1_n_581);
  ATT1_g13576 : OAI22D0BWP7T port map(A1 => ATT1_n_516, A2 => ATT1_n_450, B1 => ATT1_n_332, B2 => ATT1_n_498, ZN => ATT1_n_580);
  ATT1_g13577 : AOI22D0BWP7T port map(A1 => ATT1_n_364, A2 => ATT1_n_488, B1 => ATT1_n_532, B2 => ATT1_n_469, ZN => ATT1_n_579);
  ATT1_g13578 : MOAI22D0BWP7T port map(A1 => ATT1_n_381, A2 => ATT1_n_510, B1 => ATT1_n_478, B2 => ATT1_n_501, ZN => ATT1_n_578);
  ATT1_g13579 : MAOI22D0BWP7T port map(A1 => ATT1_n_485, A2 => ATT1_n_534, B1 => ATT1_n_408, B2 => ATT1_n_496, ZN => ATT1_n_577);
  ATT1_g13580 : MOAI22D0BWP7T port map(A1 => ATT1_n_483, A2 => ATT1_n_490, B1 => ATT1_n_514, B2 => ATT1_n_492, ZN => ATT1_n_576);
  ATT1_g13581 : AOI22D0BWP7T port map(A1 => ATT1_n_378, A2 => ATT1_n_509, B1 => ATT1_n_401, B2 => ATT1_n_491, ZN => ATT1_n_575);
  ATT1_g13582 : MOAI22D0BWP7T port map(A1 => ATT1_n_418, A2 => ATT1_n_468, B1 => ATT1_n_360, B2 => ATT1_n_522, ZN => ATT1_n_574);
  ATT1_g13583 : OAI22D0BWP7T port map(A1 => ATT1_n_406, A2 => ATT1_n_521, B1 => ATT1_n_407, B2 => ATT1_n_450, ZN => ATT1_n_573);
  ATT1_g13584 : MOAI22D0BWP7T port map(A1 => ATT1_n_454, A2 => ATT1_n_493, B1 => ATT1_n_532, B2 => ATT1_n_479, ZN => ATT1_n_572);
  ATT1_g13585 : OAI22D0BWP7T port map(A1 => ATT1_n_536, A2 => ATT1_n_466, B1 => ATT1_n_414, B2 => ATT1_n_521, ZN => ATT1_n_571);
  ATT1_g13586 : AO22D0BWP7T port map(A1 => ATT1_n_519, A2 => ATT1_n_525, B1 => ATT1_n_479, B2 => ATT1_n_387, Z => ATT1_n_570);
  ATT1_g13587 : OA22D0BWP7T port map(A1 => ATT1_n_538, A2 => ATT1_n_481, B1 => ATT1_n_489, B2 => ATT1_n_517, Z => ATT1_n_569);
  ATT1_g13588 : OAI22D0BWP7T port map(A1 => ATT1_n_515, A2 => ATT1_n_495, B1 => ATT1_n_422, B2 => ATT1_n_438, ZN => ATT1_n_568);
  ATT1_g13589 : OAI22D0BWP7T port map(A1 => ATT1_n_419, A2 => ATT1_n_521, B1 => ATT1_n_378, B2 => ATT1_n_498, ZN => ATT1_n_567);
  ATT1_g13590 : AO22D0BWP7T port map(A1 => ATT1_n_361, A2 => ATT1_n_524, B1 => ATT1_n_479, B2 => ATT1_n_405, Z => ATT1_n_566);
  ATT1_g13591 : AOI22D0BWP7T port map(A1 => ATT1_n_355, A2 => ATT1_n_39, B1 => ATT1_n_403, B2 => ATT1_n_467, ZN => ATT1_n_565);
  ATT1_g13592 : OAI22D0BWP7T port map(A1 => ATT1_n_463, A2 => ATT1_n_523, B1 => ATT1_n_332, B2 => ATT1_n_495, ZN => ATT1_n_564);
  ATT1_g13593 : OA222D0BWP7T port map(A1 => ATT1_n_515, A2 => ATT1_n_498, B1 => ATT1_n_471, B2 => ATT1_n_422, C1 => ATT1_n_450, C2 => ATT1_n_396, Z => ATT1_n_563);
  ATT1_g13594 : OA33D0BWP7T port map(A1 => ATT1_n_502, A2 => ATT1_n_429, A3 => ATT1_n_453, B1 => ATT1_n_476, B2 => ATT1_n_348, B3 => ATT1_n_384, Z => ATT1_n_586);
  ATT1_g13595 : INVD1BWP7T port map(I => ATT1_n_557, ZN => ATT1_n_556);
  ATT1_g13596 : AOI21D0BWP7T port map(A1 => ATT1_n_477, A2 => ATT1_n_390, B => ATT1_n_440, ZN => ATT1_n_554);
  ATT1_g13597 : ND4D0BWP7T port map(A1 => ATT1_n_341, A2 => ATT1_n_340, A3 => ATT1_n_468, A4 => ATT1_n_827, ZN => ATT1_n_553);
  ATT1_g13598 : NR3D0BWP7T port map(A1 => ATT1_n_478, A2 => ATT1_n_484, A3 => ATT1_n_500, ZN => ATT1_n_552);
  ATT1_g13599 : ND2D1BWP7T port map(A1 => ATT1_n_530, A2 => ATT1_n_377, ZN => ATT1_n_562);
  ATT1_g13600 : NR2XD0BWP7T port map(A1 => ATT1_n_528, A2 => ATT1_n_492, ZN => ATT1_n_561);
  ATT1_g13601 : INR2XD0BWP7T port map(A1 => ATT1_n_438, B1 => ATT1_n_528, ZN => ATT1_n_560);
  ATT1_g13602 : NR2XD0BWP7T port map(A1 => ATT1_n_499, A2 => ATT1_n_39, ZN => ATT1_n_559);
  ATT1_g13603 : NR2XD0BWP7T port map(A1 => ATT1_n_509, A2 => ATT1_n_494, ZN => ATT1_n_558);
  ATT1_g13604 : ND4D0BWP7T port map(A1 => ATT1_n_362, A2 => ATT1_n_346, A3 => ATT1_n_345, A4 => ATT1_n_464, ZN => ATT1_n_557);
  ATT1_g13605 : ND4D0BWP7T port map(A1 => ATT1_n_362, A2 => ATT1_n_346, A3 => ATT1_n_345, A4 => ATT1_n_465, ZN => ATT1_n_555);
  ATT1_g13606 : INVD0BWP7T port map(I => ATT1_n_549, ZN => ATT1_n_550);
  ATT1_g13607 : NR3D0BWP7T port map(A1 => ATT1_n_422, A2 => ATT1_n_382, A3 => ATT1_n_495, ZN => ATT1_n_548);
  ATT1_g13608 : OAI21D0BWP7T port map(A1 => ATT1_n_402, A2 => ATT1_n_368, B => ATT1_n_522, ZN => ATT1_n_547);
  ATT1_g13609 : OAI22D0BWP7T port map(A1 => ATT1_n_463, A2 => ATT1_n_496, B1 => ATT1_n_455, B2 => ATT1_n_481, ZN => ATT1_n_546);
  ATT1_g13610 : AOI21D0BWP7T port map(A1 => ATT1_n_419, A2 => ATT1_n_381, B => ATT1_n_527, ZN => ATT1_n_545);
  ATT1_g13611 : OAI21D0BWP7T port map(A1 => ATT1_n_399, A2 => ATT1_n_360, B => ATT1_n_528, ZN => ATT1_n_544);
  ATT1_g13612 : IND3D0BWP7T port map(A1 => ATT1_n_422, B1 => ATT1_n_499, B2 => ATT1_n_381, ZN => ATT1_n_543);
  ATT1_g13613 : OAI22D0BWP7T port map(A1 => ATT1_n_477, A2 => ATT1_n_468, B1 => ATT1_n_483, B2 => ATT1_n_466, ZN => ATT1_n_542);
  ATT1_g13614 : MAOI22D0BWP7T port map(A1 => ATT1_n_394, A2 => ATT1_n_491, B1 => ATT1_n_418, B2 => ATT1_n_500, ZN => ATT1_n_541);
  ATT1_g13615 : AO22D0BWP7T port map(A1 => ATT1_n_361, A2 => ATT1_n_497, B1 => ATT1_n_451, B2 => ATT1_n_405, Z => ATT1_n_540);
  ATT1_g13616 : NR4D0BWP7T port map(A1 => ATT1_n_478, A2 => ATT1_n_392, A3 => ATT1_n_350, A4 => FE_OFN2_ATT1_n_301, ZN => ATT1_n_551);
  ATT1_g13617 : NR3D0BWP7T port map(A1 => ATT1_n_453, A2 => ATT1_n_429, A3 => ATT1_n_40, ZN => ATT1_n_549);
  ATT1_g13618 : CKND1BWP7T port map(I => ATT1_n_535, ZN => ATT1_n_536);
  ATT1_g13619 : INVD0BWP7T port map(I => ATT1_n_530, ZN => ATT1_n_529);
  ATT1_g13620 : INVD0BWP7T port map(I => ATT1_n_528, ZN => ATT1_n_527);
  ATT1_g13621 : INVD1BWP7T port map(I => ATT1_n_525, ZN => ATT1_n_526);
  ATT1_g13622 : INVD1BWP7T port map(I => ATT1_n_524, ZN => ATT1_n_523);
  ATT1_g13623 : INVD1BWP7T port map(I => ATT1_n_522, ZN => ATT1_n_521);
  ATT1_g13624 : ND2D0BWP7T port map(A1 => ATT1_n_477, A2 => ATT1_n_426, ZN => ATT1_n_520);
  ATT1_g13625 : NR2XD0BWP7T port map(A1 => ATT1_n_488, A2 => ATT1_n_469, ZN => ATT1_n_539);
  ATT1_g13626 : NR4D0BWP7T port map(A1 => ATT1_n_478, A2 => ATT1_n_398, A3 => ATT1_n_389, A4 => ATT1_n_337, ZN => ATT1_n_538);
  ATT1_g13627 : NR4D0BWP7T port map(A1 => ATT1_n_478, A2 => ATT1_n_411, A3 => ATT1_n_343, A4 => ATT1_n_337, ZN => ATT1_n_537);
  ATT1_g13628 : ND2D1BWP7T port map(A1 => ATT1_n_477, A2 => ATT1_n_414, ZN => ATT1_n_535);
  ATT1_g13629 : ND2D1BWP7T port map(A1 => ATT1_n_481, A2 => ATT1_n_489, ZN => ATT1_n_534);
  ATT1_g13630 : NR2XD0BWP7T port map(A1 => ATT1_n_492, A2 => ATT1_n_501, ZN => ATT1_n_533);
  ATT1_g13631 : NR2D1BWP7T port map(A1 => ATT1_n_484, A2 => ATT1_n_360, ZN => ATT1_n_532);
  ATT1_g13632 : NR2XD0BWP7T port map(A1 => ATT1_n_492, A2 => ATT1_n_430, ZN => ATT1_n_531);
  ATT1_g13633 : NR2D1BWP7T port map(A1 => ATT1_n_478, A2 => ATT1_n_383, ZN => ATT1_n_530);
  ATT1_g13634 : IND2D1BWP7T port map(A1 => ATT1_n_430, B1 => ATT1_n_40, ZN => ATT1_n_528);
  ATT1_g13635 : ND2D1BWP7T port map(A1 => ATT1_n_490, A2 => ATT1_n_441, ZN => ATT1_n_525);
  ATT1_g13636 : ND2D1BWP7T port map(A1 => ATT1_n_500, A2 => ATT1_n_438, ZN => ATT1_n_524);
  ATT1_g13637 : ND2D1BWP7T port map(A1 => ATT1_n_502, A2 => ATT1_n_444, ZN => ATT1_n_522);
  ATT1_g13638 : INVD0BWP7T port map(I => ATT1_n_518, ZN => diry2new1(7));
  ATT1_g13639 : INVD0BWP7T port map(I => ATT1_n_512, ZN => ATT1_n_511);
  ATT1_g13640 : INVD1BWP7T port map(I => ATT1_n_510, ZN => ATT1_n_509);
  ATT1_g13641 : INVD1BWP7T port map(I => ATT1_n_39, ZN => ATT1_n_508);
  ATT1_g13642 : ND3D0BWP7T port map(A1 => ATT1_n_452, A2 => ATT1_n_313, A3 => ATT1_n_309, ZN => ATT1_n_507);
  ATT1_g13643 : MOAI22D0BWP7T port map(A1 => ATT1_n_422, A2 => ATT1_n_442, B1 => ATT1_n_401, B2 => ATT1_n_467, ZN => ATT1_n_506);
  ATT1_g13644 : OAI22D0BWP7T port map(A1 => ATT1_n_454, A2 => ATT1_n_438, B1 => ATT1_n_443, B2 => ATT1_n_441, ZN => ATT1_n_505);
  ATT1_g13645 : OAI22D0BWP7T port map(A1 => ATT1_n_454, A2 => ATT1_n_440, B1 => ATT1_n_443, B2 => ATT1_n_442, ZN => ATT1_n_504);
  ATT1_g13646 : AO21D0BWP7T port map(A1 => ATT1_n_421, A2 => ATT1_n_379, B => ATT1_n_40, Z => ATT1_n_503);
  ATT1_g13647 : ND4D0BWP7T port map(A1 => ATT1_n_452, A2 => ATT1_n_388, A3 => ATT1_n_393, A4 => ATT1_n_344, ZN => ATT1_n_519);
  ATT1_g13648 : ND3D0BWP7T port map(A1 => ATT1_n_316, A2 => ATT1_n_320, A3 => ATT1_n_817, ZN => ATT1_n_518);
  ATT1_g13649 : ND4D0BWP7T port map(A1 => ATT1_n_432, A2 => ATT1_n_344, A3 => ATT1_n_349, A4 => ATT1_n_300, ZN => ATT1_n_517);
  ATT1_g13650 : ND4D0BWP7T port map(A1 => ATT1_n_432, A2 => ATT1_n_393, A3 => ATT1_n_309, A4 => ATT1_n_300, ZN => ATT1_n_516);
  ATT1_g13651 : NR3D0BWP7T port map(A1 => ATT1_n_478, A2 => ATT1_n_403, A3 => ATT1_n_382, ZN => ATT1_n_515);
  ATT1_g13652 : ND4D0BWP7T port map(A1 => ATT1_n_452, A2 => ATT1_n_375, A3 => ATT1_n_370, A4 => ATT1_n_319, ZN => ATT1_n_514);
  ATT1_g13653 : AOI21D0BWP7T port map(A1 => ATT1_n_474, A2 => ATT1_n_444, B => ATT1_n_336, ZN => ATT1_n_513);
  ATT1_g13654 : ND3D0BWP7T port map(A1 => ATT1_n_477, A2 => ATT1_n_427, A3 => ATT1_n_381, ZN => ATT1_n_512);
  ATT1_g13655 : ND3D0BWP7T port map(A1 => ATT1_n_316, A2 => ATT1_n_326, A3 => ATT1_n_470, ZN => ATT1_n_510);
  ATT1_g13657 : INVD1BWP7T port map(I => ATT1_n_501, ZN => ATT1_n_500);
  ATT1_g13658 : INVD1BWP7T port map(I => ATT1_n_499, ZN => ATT1_n_498);
  ATT1_g13659 : INVD1BWP7T port map(I => ATT1_n_497, ZN => ATT1_n_496);
  ATT1_g13660 : INVD1BWP7T port map(I => ATT1_n_495, ZN => ATT1_n_494);
  ATT1_g13661 : INVD1BWP7T port map(I => ATT1_n_493, ZN => ATT1_n_492);
  ATT1_g13662 : INVD1BWP7T port map(I => ATT1_n_491, ZN => ATT1_n_490);
  ATT1_g13663 : INVD1BWP7T port map(I => ATT1_n_489, ZN => ATT1_n_488);
  ATT1_g13664 : IND2D1BWP7T port map(A1 => ATT1_n_474, B1 => ATT1_n_336, ZN => ATT1_n_502);
  ATT1_g13665 : NR2D1BWP7T port map(A1 => ATT1_n_266, A2 => ATT1_n_475, ZN => ATT1_n_501);
  ATT1_g13666 : NR2D1BWP7T port map(A1 => ATT1_n_341, A2 => ATT1_n_473, ZN => ATT1_n_499);
  ATT1_g13667 : ND2D1BWP7T port map(A1 => ATT1_n_468, A2 => ATT1_n_440, ZN => ATT1_n_497);
  ATT1_g13668 : IND2D1BWP7T port map(A1 => ATT1_n_341, B1 => ATT1_n_470, ZN => ATT1_n_495);
  ATT1_g13669 : IND2D1BWP7T port map(A1 => ATT1_n_340, B1 => ATT1_n_817, ZN => ATT1_n_493);
  ATT1_g13670 : NR2D1BWP7T port map(A1 => ATT1_n_267, A2 => ATT1_n_475, ZN => ATT1_n_491);
  ATT1_g13671 : IND2D1BWP7T port map(A1 => ATT1_n_340, B1 => ATT1_n_827, ZN => ATT1_n_489);
  ATT1_g13672 : CKND1BWP7T port map(I => ATT1_n_485, ZN => ATT1_n_486);
  ATT1_g13673 : INVD1BWP7T port map(I => ATT1_n_482, ZN => ATT1_n_481);
  ATT1_g13674 : INVD1BWP7T port map(I => ATT1_n_480, ZN => ATT1_n_479);
  ATT1_g13675 : INVD1BWP7T port map(I => ATT1_n_478, ZN => ATT1_n_477);
  ATT1_g13676 : IND3D1BWP7T port map(A1 => ATT1_n_444, B1 => ATT1_n_353, B2 => ATT1_n_424, ZN => ATT1_n_476);
  ATT1_g13677 : NR2D1BWP7T port map(A1 => ATT1_n_336, A2 => ATT1_n_457, ZN => ATT1_n_487);
  ATT1_g13678 : ND2D1BWP7T port map(A1 => ATT1_n_452, A2 => ATT1_n_433, ZN => ATT1_n_485);
  ATT1_g13679 : ND3D0BWP7T port map(A1 => ATT1_n_428, A2 => ATT1_n_322, A3 => ATT1_n_324, ZN => ATT1_n_484);
  ATT1_g13680 : IND2D1BWP7T port map(A1 => ATT1_n_456, B1 => ATT1_n_313, ZN => ATT1_n_483);
  ATT1_g13682 : ND2D1BWP7T port map(A1 => ATT1_n_466, A2 => ATT1_n_442, ZN => ATT1_n_482);
  ATT1_g13683 : ND3D0BWP7T port map(A1 => ATT1_n_302, A2 => ATT1_n_285, A3 => ATT1_n_423, ZN => ATT1_n_480);
  ATT1_g13684 : ND2D1BWP7T port map(A1 => ATT1_n_452, A2 => ATT1_n_336, ZN => ATT1_n_478);
  ATT1_g13685 : INVD1BWP7T port map(I => ATT1_n_469, ZN => ATT1_n_468);
  ATT1_g13686 : INVD1BWP7T port map(I => ATT1_n_467, ZN => ATT1_n_466);
  ATT1_g13687 : NR2XD0BWP7T port map(A1 => ATT1_n_371, A2 => ATT1_n_449, ZN => ATT1_n_465);
  ATT1_g13688 : NR2XD0BWP7T port map(A1 => ATT1_n_371, A2 => ATT1_n_446, ZN => ATT1_n_464);
  ATT1_g13689 : CKND2D1BWP7T port map(A1 => ATT1_n_307, A2 => ATT1_n_423, ZN => ATT1_n_475);
  ATT1_g13690 : ND2D1BWP7T port map(A1 => ATT1_n_363, A2 => ATT1_n_425, ZN => ATT1_n_474);
  ATT1_g13691 : NR2D1BWP7T port map(A1 => ATT1_n_425, A2 => ATT1_n_412, ZN => ATT1_n_473);
  ATT1_g13692 : IND2D1BWP7T port map(A1 => ATT1_n_441, B1 => ATT1_n_361, ZN => ATT1_n_472);
  ATT1_g13693 : CKAN2D1BWP7T port map(A1 => ATT1_n_440, A2 => ATT1_n_442, Z => ATT1_n_471);
  ATT1_g13694 : OR2D1BWP7T port map(A1 => ATT1_n_423, A2 => ATT1_n_413, Z => ATT1_n_470);
  ATT1_g13695 : CKND2D1BWP7T port map(A1 => ATT1_n_404, A2 => ATT1_n_446, ZN => ATT1_n_827);
  ATT1_g13696 : IND2D1BWP7T port map(A1 => ATT1_n_423, B1 => ATT1_n_449, ZN => ATT1_n_817);
  ATT1_g13697 : NR2XD0BWP7T port map(A1 => ATT1_n_266, A2 => ATT1_n_448, ZN => ATT1_n_469);
  ATT1_g13698 : NR2XD0BWP7T port map(A1 => ATT1_n_267, A2 => ATT1_n_448, ZN => ATT1_n_467);
  ATT1_g13700 : INVD1BWP7T port map(I => ATT1_n_454, ZN => ATT1_n_453);
  ATT1_g13701 : INVD1BWP7T port map(I => ATT1_n_451, ZN => ATT1_n_450);
  ATT1_g13702 : IND4D0BWP7T port map(A1 => ATT1_n_389, B1 => ATT1_n_338, B2 => ATT1_n_365, B3 => ATT1_n_393, ZN => ATT1_n_463);
  ATT1_g13703 : NR2D0BWP7T port map(A1 => ATT1_n_429, A2 => ATT1_n_355, ZN => ATT1_n_462);
  ATT1_g13704 : CKAN2D1BWP7T port map(A1 => ATT1_n_427, A2 => ATT1_n_377, Z => ATT1_n_461);
  ATT1_g13705 : CKAN2D1BWP7T port map(A1 => ATT1_n_427, A2 => ATT1_n_400, Z => ATT1_n_460);
  ATT1_g13706 : IND4D0BWP7T port map(A1 => ATT1_n_373, B1 => ATT1_n_300, B2 => ATT1_n_370, B3 => ATT1_n_393, ZN => ATT1_n_459);
  ATT1_g13707 : IND2D1BWP7T port map(A1 => ATT1_n_442, B1 => ATT1_n_361, ZN => ATT1_n_458);
  ATT1_g13708 : IND3D1BWP7T port map(A1 => ATT1_n_371, B1 => ATT1_n_423, B2 => ATT1_n_305, ZN => ATT1_n_457);
  ATT1_g13709 : ND2D1BWP7T port map(A1 => ATT1_n_428, A2 => ATT1_n_375, ZN => ATT1_n_456);
  ATT1_g13710 : ND2D1BWP7T port map(A1 => ATT1_n_428, A2 => ATT1_n_370, ZN => ATT1_n_455);
  ATT1_g13711 : NR3D0BWP7T port map(A1 => ATT1_n_402, A2 => ATT1_n_343, A3 => ATT1_n_350, ZN => ATT1_n_454);
  ATT1_g13712 : IND2D1BWP7T port map(A1 => ATT1_n_417, B1 => ATT1_n_424, ZN => ATT1_n_452);
  ATT1_g13713 : INR3D0BWP7T port map(A1 => ATT1_n_285, B1 => ATT1_n_404, B2 => ATT1_n_295, ZN => ATT1_n_451);
  ATT1_g13714 : INVD0BWP7T port map(I => ATT1_n_440, ZN => ATT1_n_439);
  ATT1_g13715 : INR2XD0BWP7T port map(A1 => ATT1_n_421, B1 => ATT1_n_368, ZN => ATT1_n_437);
  ATT1_g13716 : CKAN2D1BWP7T port map(A1 => ATT1_n_406, A2 => ATT1_n_381, Z => ATT1_n_436);
  ATT1_g13717 : ND2D1BWP7T port map(A1 => ATT1_n_347, A2 => ATT1_n_413, ZN => ATT1_n_449);
  ATT1_g13718 : IND2D1BWP7T port map(A1 => ATT1_n_404, B1 => ATT1_n_307, ZN => ATT1_n_448);
  ATT1_g13719 : NR2XD0BWP7T port map(A1 => ATT1_n_401, A2 => ATT1_n_382, ZN => ATT1_n_447);
  ATT1_g13720 : ND2D1BWP7T port map(A1 => ATT1_n_347, A2 => ATT1_n_412, ZN => ATT1_n_446);
  ATT1_g13721 : CKAN2D1BWP7T port map(A1 => ATT1_n_415, A2 => ATT1_n_381, Z => ATT1_n_445);
  ATT1_g13722 : IND2D1BWP7T port map(A1 => ATT1_n_345, B1 => ATT1_n_412, ZN => ATT1_n_444);
  ATT1_g13723 : CKAN2D1BWP7T port map(A1 => ATT1_n_416, A2 => ATT1_n_313, Z => ATT1_n_443);
  ATT1_g13724 : IND2D1BWP7T port map(A1 => ATT1_n_346, B1 => ATT1_n_412, ZN => ATT1_n_442);
  ATT1_g13725 : IND2D1BWP7T port map(A1 => ATT1_n_346, B1 => ATT1_n_413, ZN => ATT1_n_441);
  ATT1_g13726 : IND2D1BWP7T port map(A1 => ATT1_n_362, B1 => ATT1_n_412, ZN => ATT1_n_440);
  ATT1_g13727 : IND2D1BWP7T port map(A1 => ATT1_n_362, B1 => ATT1_n_413, ZN => ATT1_n_438);
  ATT1_g13728 : INR2XD0BWP7T port map(A1 => ATT1_n_393, B1 => ATT1_n_402, ZN => ATT1_n_435);
  ATT1_g13729 : NR2XD0BWP7T port map(A1 => ATT1_n_399, A2 => ATT1_n_383, ZN => ATT1_n_434);
  ATT1_g13730 : INR2XD0BWP7T port map(A1 => ATT1_n_379, B1 => ATT1_n_402, ZN => ATT1_n_433);
  ATT1_g13731 : NR3D0BWP7T port map(A1 => ATT1_n_395, A2 => ATT1_n_335, A3 => ATT1_n_337, ZN => ATT1_n_432);
  ATT1_g13732 : NR2XD0BWP7T port map(A1 => ATT1_n_399, A2 => ATT1_n_403, ZN => ATT1_n_431);
  ATT1_g13733 : INR2D1BWP7T port map(A1 => ATT1_n_413, B1 => ATT1_n_345, ZN => ATT1_n_430);
  ATT1_g13734 : ND2D1BWP7T port map(A1 => ATT1_n_400, A2 => ATT1_n_300, ZN => ATT1_n_429);
  ATT1_g13735 : NR3D0BWP7T port map(A1 => ATT1_n_392, A2 => ATT1_n_373, A3 => FE_OFN2_ATT1_n_301, ZN => ATT1_n_428);
  ATT1_g13736 : NR2XD0BWP7T port map(A1 => ATT1_n_401, A2 => ATT1_n_360, ZN => ATT1_n_427);
  ATT1_g13737 : NR4D0BWP7T port map(A1 => ATT1_n_389, A2 => ATT1_n_343, A3 => ATT1_n_351, A4 => ATT1_n_348, ZN => ATT1_n_426);
  ATT1_g13738 : INR3D0BWP7T port map(A1 => ATT1_n_305, B1 => ATT1_n_404, B2 => ATT1_n_339, ZN => ATT1_n_425);
  ATT1_g13739 : NR2XD0BWP7T port map(A1 => ATT1_n_402, A2 => ATT1_n_392, ZN => ATT1_n_424);
  ATT1_g13740 : NR3D0BWP7T port map(A1 => ATT1_n_358, A2 => ATT1_n_386, A3 => orientationp1, ZN => ATT1_n_423);
  ATT1_g13741 : OR2D1BWP7T port map(A1 => ATT1_n_401, A2 => FE_OFN2_ATT1_n_301, Z => ATT1_n_422);
  ATT1_g13742 : OR2D1BWP7T port map(A1 => ATT1_n_392, A2 => ATT1_n_395, Z => ATT1_n_411);
  ATT1_g13743 : INR2XD0BWP7T port map(A1 => ATT1_n_319, B1 => ATT1_n_395, ZN => ATT1_n_421);
  ATT1_g13744 : INR2XD0BWP7T port map(A1 => ATT1_n_322, B1 => ATT1_n_389, ZN => ATT1_n_420);
  ATT1_g13745 : NR2XD0BWP7T port map(A1 => ATT1_n_391, A2 => ATT1_n_355, ZN => ATT1_n_419);
  ATT1_g13746 : NR2XD0BWP7T port map(A1 => ATT1_n_394, A2 => ATT1_n_383, ZN => ATT1_n_418);
  ATT1_g13747 : IND2D1BWP7T port map(A1 => ATT1_n_384, B1 => ATT1_n_322, ZN => ATT1_n_417);
  ATT1_g13748 : NR2XD0BWP7T port map(A1 => ATT1_n_389, A2 => ATT1_n_392, ZN => ATT1_n_416);
  ATT1_g13749 : NR2XD0BWP7T port map(A1 => ATT1_n_383, A2 => ATT1_n_355, ZN => ATT1_n_415);
  ATT1_g13750 : NR2XD0BWP7T port map(A1 => ATT1_n_391, A2 => ATT1_n_378, ZN => ATT1_n_414);
  ATT1_g13751 : INR2XD0BWP7T port map(A1 => orientationp1, B1 => ATT1_n_386, ZN => ATT1_n_413);
  ATT1_g13752 : NR2XD0BWP7T port map(A1 => ATT1_n_385, A2 => orientationp2, ZN => ATT1_n_412);
  ATT1_g13753 : INVD1BWP7T port map(I => ATT1_n_400, ZN => ATT1_n_399);
  ATT1_g13754 : ND2D1BWP7T port map(A1 => ATT1_n_393, A2 => ATT1_n_318, ZN => ATT1_n_398);
  ATT1_g13755 : IND2D1BWP7T port map(A1 => ATT1_n_384, B1 => ATT1_n_379, ZN => ATT1_n_410);
  ATT1_g13756 : NR2XD0BWP7T port map(A1 => ATT1_n_389, A2 => ATT1_n_368, ZN => ATT1_n_409);
  ATT1_g13757 : OR2D1BWP7T port map(A1 => ATT1_n_384, A2 => ATT1_n_392, Z => ATT1_n_408);
  ATT1_g13758 : IND4D0BWP7T port map(A1 => ATT1_n_310, B1 => ATT1_n_332, B2 => ATT1_n_334, B3 => ATT1_n_365, ZN => ATT1_n_407);
  ATT1_g13759 : INR2XD0BWP7T port map(A1 => ATT1_n_388, B1 => ATT1_n_368, ZN => ATT1_n_406);
  ATT1_g13760 : NR2D1BWP7T port map(A1 => ATT1_n_382, A2 => FE_OFN2_ATT1_n_301, ZN => ATT1_n_405);
  ATT1_g13761 : IND3D1BWP7T port map(A1 => ATT1_n_385, B1 => orientationp2, B2 => ATT1_n_357, ZN => ATT1_n_404);
  ATT1_g13762 : OR3D1BWP7T port map(A1 => ATT1_n_310, A2 => ATT1_n_350, A3 => ATT1_n_389, Z => ATT1_n_403);
  ATT1_g13763 : IND2D1BWP7T port map(A1 => ATT1_n_389, B1 => ATT1_n_319, ZN => ATT1_n_402);
  ATT1_g13764 : OR2D1BWP7T port map(A1 => ATT1_n_389, A2 => ATT1_n_333, Z => ATT1_n_401);
  ATT1_g13765 : NR2XD0BWP7T port map(A1 => ATT1_n_382, A2 => ATT1_n_378, ZN => ATT1_n_400);
  ATT1_g13766 : INVD0BWP7T port map(I => ATT1_n_396, ZN => ATT1_n_397);
  ATT1_g13767 : INVD0BWP7T port map(I => ATT1_n_391, ZN => ATT1_n_390);
  ATT1_g13768 : NR2XD0BWP7T port map(A1 => ATT1_n_378, A2 => ATT1_n_355, ZN => ATT1_n_396);
  ATT1_g13769 : ND2D1BWP7T port map(A1 => ATT1_n_375, A2 => ATT1_n_324, ZN => ATT1_n_395);
  ATT1_g13770 : IND2D1BWP7T port map(A1 => ATT1_n_351, B1 => ATT1_n_377, ZN => ATT1_n_394);
  ATT1_g13771 : AN2D1BWP7T port map(A1 => ATT1_n_376, A2 => ATT1_n_349, Z => ATT1_n_393);
  ATT1_g13772 : ND2D1BWP7T port map(A1 => ATT1_n_376, A2 => ATT1_n_369, ZN => ATT1_n_392);
  ATT1_g13773 : ND2D1BWP7T port map(A1 => ATT1_n_375, A2 => ATT1_n_318, ZN => ATT1_n_391);
  ATT1_g13774 : OR2D1BWP7T port map(A1 => ATT1_n_373, A2 => ATT1_n_374, Z => ATT1_n_389);
  ATT1_g13775 : INVD1BWP7T port map(I => ATT1_n_382, ZN => ATT1_n_381);
  ATT1_g13776 : AN3D1BWP7T port map(A1 => ATT1_n_372, A2 => ATT1_n_318, A3 => ATT1_n_319, Z => ATT1_n_388);
  ATT1_g13777 : IND4D0BWP7T port map(A1 => ATT1_n_373, B1 => ATT1_n_309, B2 => ATT1_n_322, B3 => ATT1_n_359, ZN => ATT1_n_387);
  ATT1_g13778 : OAI21D0BWP7T port map(A1 => ATT1_at1a, A2 => ATT1_at1b, B => ATT1_n_380, ZN => ATT1_n_386);
  ATT1_g13779 : OAI21D0BWP7T port map(A1 => ATT1_at2a, A2 => ATT1_at2b, B => ATT1_n_380, ZN => ATT1_n_385);
  ATT1_g13780 : ND3D0BWP7T port map(A1 => ATT1_n_370, A2 => ATT1_n_324, A3 => ATT1_n_300, ZN => ATT1_n_384);
  ATT1_g13781 : IND2D1BWP7T port map(A1 => ATT1_n_373, B1 => ATT1_n_324, ZN => ATT1_n_383);
  ATT1_g13782 : ND2D1BWP7T port map(A1 => ATT1_n_376, A2 => ATT1_n_332, ZN => ATT1_n_382);
  ATT1_g13783 : INVD1BWP7T port map(I => ATT1_n_378, ZN => ATT1_n_377);
  ATT1_g13784 : AO211D0BWP7T port map(A1 => ATT1_n_320, A2 => ATT1_n_304, B => ATT1_n_356, C => ATT1_n_354, Z => ATT1_n_380);
  ATT1_g13785 : NR2XD0BWP7T port map(A1 => ATT1_n_368, A2 => ATT1_n_331, ZN => ATT1_n_379);
  ATT1_g13786 : ND2D1BWP7T port map(A1 => ATT1_n_369, A2 => ATT1_n_349, ZN => ATT1_n_378);
  ATT1_g13787 : INVD1BWP7T port map(I => ATT1_n_375, ZN => ATT1_n_374);
  ATT1_g13788 : INVD1BWP7T port map(I => ATT1_n_372, ZN => ATT1_n_373);
  ATT1_g13789 : ND3D0BWP7T port map(A1 => ATT1_n_356, A2 => ATT1_n_300, A3 => ATT1_n_288, ZN => ATT1_n_376);
  ATT1_g13790 : ND3D0BWP7T port map(A1 => ATT1_n_356, A2 => ATT1_n_278, A3 => ATT1_n_233, ZN => ATT1_n_375);
  ATT1_g13791 : ND3D0BWP7T port map(A1 => ATT1_n_356, A2 => ATT1_n_278, A3 => ATT1_n_232, ZN => ATT1_n_372);
  ATT1_g13792 : INVD1BWP7T port map(I => ATT1_n_369, ZN => ATT1_n_368);
  ATT1_g13793 : ND2D1BWP7T port map(A1 => ATT1_n_363, A2 => ATT1_n_340, ZN => ATT1_n_371);
  ATT1_g13794 : AN2D1BWP7T port map(A1 => ATT1_n_359, A2 => ATT1_n_344, Z => ATT1_n_370);
  ATT1_g13795 : ND2D1BWP7T port map(A1 => ATT1_n_356, A2 => ATT1_n_289, ZN => ATT1_n_369);
  ATT1_g13796 : INVD0BWP7T port map(I => ATT1_n_366, ZN => ATT1_n_367);
  ATT1_g13798 : IND3D1BWP7T port map(A1 => ATT1_n_351, B1 => ATT1_n_322, B2 => ATT1_n_324, ZN => ATT1_n_366);
  ATT1_g13799 : NR3D0BWP7T port map(A1 => ATT1_n_343, A2 => ATT1_n_335, A3 => FE_OFN2_ATT1_n_301, ZN => ATT1_n_365);
  ATT1_g13800 : NR2D1BWP7T port map(A1 => ATT1_n_360, A2 => FE_OFN2_ATT1_n_301, ZN => ATT1_n_364);
  ATT1_g13801 : NR2XD0BWP7T port map(A1 => ATT1_n_352, A2 => ATT1_n_326, ZN => ATT1_n_363);
  ATT1_g13802 : AOI21D0BWP7T port map(A1 => ATT1_n_325, A2 => ATT1_n_198, B => ATT1_n_342, ZN => ATT1_n_362);
  ATT1_g13803 : NR2D1BWP7T port map(A1 => ATT1_n_351, A2 => FE_OFN2_ATT1_n_301, ZN => ATT1_n_361);
  ATT1_g13804 : ND2D1BWP7T port map(A1 => ATT1_n_344, A2 => ATT1_n_309, ZN => ATT1_n_360);
  ATT1_g13805 : INVD0BWP7T port map(I => ATT1_n_357, ZN => ATT1_n_358);
  ATT1_g13806 : AOI211XD0BWP7T port map(A1 => ATT1_n_278, A2 => ATT1_n_250, B => ATT1_n_328, C => ATT1_n_304, ZN => ATT1_n_354);
  ATT1_g13807 : AN3D0BWP7T port map(A1 => ATT1_n_336, A2 => ATT1_n_338, A3 => ATT1_n_318, Z => ATT1_n_359);
  ATT1_g13808 : OAI22D0BWP7T port map(A1 => ATT1_n_330, A2 => ATT1_n_296, B1 => ATT1_n_314, B2 => ATT1_n_264, ZN => ATT1_n_357);
  ATT1_g13809 : NR3D0BWP7T port map(A1 => ATT1_n_329, A2 => ATT1_n_304, A3 => ATT1_n_284, ZN => ATT1_n_356);
  ATT1_g13810 : ND3D0BWP7T port map(A1 => ATT1_n_344, A2 => ATT1_n_338, A3 => ATT1_n_319, ZN => ATT1_n_355);
  ATT1_g13811 : INVD0BWP7T port map(I => ATT1_n_349, ZN => ATT1_n_348);
  ATT1_g13812 : ND2D1BWP7T port map(A1 => ATT1_n_331, A2 => ATT1_n_161, ZN => ATT1_n_353);
  ATT1_g13813 : ND2D1BWP7T port map(A1 => ATT1_n_341, A2 => ATT1_n_316, ZN => ATT1_n_352);
  ATT1_g13814 : IND2D1BWP7T port map(A1 => ATT1_n_310, B1 => ATT1_n_338, ZN => ATT1_n_351);
  ATT1_g13815 : ND2D1BWP7T port map(A1 => ATT1_n_338, A2 => ATT1_n_334, ZN => ATT1_n_350);
  ATT1_g13816 : ND2D1BWP7T port map(A1 => ATT1_n_332, A2 => ATT1_n_323, ZN => ATT1_n_349);
  ATT1_g13817 : INVD1BWP7T port map(I => ATT1_n_344, ZN => ATT1_n_343);
  ATT1_g13818 : NR4D0BWP7T port map(A1 => ATT1_n_311, A2 => ATT1_n_291, A3 => ATT1_n_266, A4 => ATT1_n_121, ZN => ATT1_n_342);
  ATT1_g13819 : OAI211D1BWP7T port map(A1 => ATT1_n_270, A2 => ATT1_n_311, B => ATT1_n_321, C => ATT1_n_314, ZN => ATT1_n_347);
  ATT1_g13820 : IND3D1BWP7T port map(A1 => ATT1_n_198, B1 => ATT1_n_196, B2 => ATT1_n_325, ZN => ATT1_n_346);
  ATT1_g13821 : MAOI22D0BWP7T port map(A1 => ATT1_n_325, A2 => ATT1_n_195, B1 => ATT1_n_314, B2 => ATT1_n_267, ZN => ATT1_n_345);
  ATT1_g13822 : ND3D0BWP7T port map(A1 => ATT1_n_327, A2 => ATT1_n_278, A3 => ATT1_n_233, ZN => ATT1_n_344);
  ATT1_g13823 : INVD1BWP7T port map(I => ATT1_n_339, ZN => ATT1_n_340);
  ATT1_g13824 : INVD1BWP7T port map(I => ATT1_n_338, ZN => ATT1_n_337);
  ATT1_g13825 : INVD0BWP7T port map(I => ATT1_n_336, ZN => ATT1_n_335);
  ATT1_g13826 : OR2D1BWP7T port map(A1 => ATT1_n_321, A2 => ATT1_n_179, Z => ATT1_n_341);
  ATT1_g13827 : NR2D1BWP7T port map(A1 => ATT1_n_321, A2 => ATT1_n_178, ZN => ATT1_n_339);
  ATT1_g13828 : ND2D1BWP7T port map(A1 => ATT1_n_327, A2 => ATT1_n_232, ZN => ATT1_n_338);
  ATT1_g13829 : IND2D1BWP7T port map(A1 => ATT1_n_278, B1 => ATT1_n_327, ZN => ATT1_n_336);
  ATT1_g13830 : CKND1BWP7T port map(I => ATT1_n_333, ZN => ATT1_n_334);
  ATT1_g13831 : INVD1BWP7T port map(I => ATT1_n_332, ZN => ATT1_n_331);
  ATT1_g13832 : AOI31D0BWP7T port map(A1 => ATT1_n_306, A2 => ATT1_n_248, A3 => ATT1_n_178, B => ATT1_n_307, ZN => ATT1_n_330);
  ATT1_g13833 : AOI21D0BWP7T port map(A1 => ATT1_n_315, A2 => ATT1_n_110, B => ATT1_n_312, ZN => ATT1_n_329);
  ATT1_g13834 : AOI21D0BWP7T port map(A1 => ATT1_n_315, A2 => ATT1_n_78, B => ATT1_n_312, ZN => ATT1_n_328);
  ATT1_g13835 : ND2D1BWP7T port map(A1 => ATT1_n_318, A2 => ATT1_n_324, ZN => ATT1_n_333);
  ATT1_g13836 : ND2D1BWP7T port map(A1 => ATT1_n_323, A2 => ATT1_n_233, ZN => ATT1_n_332);
  ATT1_g13838 : INVD1BWP7T port map(I => ATT1_n_323, ZN => ATT1_n_322);
  ATT1_g13839 : CKAN2D1BWP7T port map(A1 => ATT1_n_304, A2 => ATT1_n_313, Z => ATT1_n_327);
  ATT1_g13840 : NR2D1BWP7T port map(A1 => ATT1_n_314, A2 => ATT1_n_266, ZN => ATT1_n_326);
  ATT1_g13841 : INR2D1BWP7T port map(A1 => ATT1_n_248, B1 => ATT1_n_314, ZN => ATT1_n_325);
  ATT1_g13842 : IND2D1BWP7T port map(A1 => ATT1_n_313, B1 => ATT1_n_289, ZN => ATT1_n_324);
  ATT1_g13843 : INR2XD0BWP7T port map(A1 => ATT1_n_278, B1 => ATT1_n_313, ZN => ATT1_n_323);
  ATT1_g13845 : INVD1BWP7T port map(I => ATT1_n_317, ZN => ATT1_n_316);
  ATT1_g13846 : IND3D1BWP7T port map(A1 => ATT1_n_296, B1 => ATT1_n_248, B2 => ATT1_n_307, ZN => ATT1_n_321);
  ATT1_g13847 : OAI31D0BWP7T port map(A1 => ATT1_n_282, A2 => ATT1_n_294, A3 => ATT1_n_303, B => ATT1_n_313, ZN => ATT1_n_320);
  ATT1_g13848 : INR2XD0BWP7T port map(A1 => ATT1_n_309, B1 => ATT1_n_310, ZN => ATT1_n_319);
  ATT1_g13849 : IND2D1BWP7T port map(A1 => ATT1_n_313, B1 => ATT1_n_288, ZN => ATT1_n_318);
  ATT1_g13850 : NR3D0BWP7T port map(A1 => ATT1_n_308, A2 => ATT1_n_266, A3 => ATT1_n_121, ZN => ATT1_n_317);
  ATT1_g13851 : AN2D0BWP7T port map(A1 => ATT1_n_303, A2 => ATT1_n_114, Z => ATT1_n_315);
  ATT1_g13852 : OR2D1BWP7T port map(A1 => ATT1_n_308, A2 => ATT1_n_302, Z => ATT1_n_314);
  ATT1_g13853 : OR2D1BWP7T port map(A1 => ATT1_n_303, A2 => ATT1_n_299, Z => ATT1_n_313);
  ATT1_g13854 : OA211D0BWP7T port map(A1 => ATT1_n_77, A2 => ATT1_n_114, B => ATT1_n_303, C => ATT1_n_286, Z => ATT1_n_312);
  ATT1_g13855 : ND4D0BWP7T port map(A1 => ATT1_n_296, A2 => ATT1_n_295, A3 => ATT1_n_279, A4 => ATT1_n_258, ZN => ATT1_n_311);
  ATT1_g13856 : AN3D1BWP7T port map(A1 => ATT1_n_303, A2 => ATT1_n_284, A3 => ATT1_n_289, Z => ATT1_n_310);
  ATT1_g13857 : ND3D0BWP7T port map(A1 => ATT1_n_303, A2 => ATT1_n_284, A3 => ATT1_n_288, ZN => ATT1_n_309);
  ATT1_g13858 : NR3D0BWP7T port map(A1 => ATT1_n_295, A2 => ATT1_n_279, A3 => ATT1_n_257, ZN => ATT1_n_306);
  ATT1_g13859 : ND2D1BWP7T port map(A1 => ATT1_n_296, A2 => ATT1_n_291, ZN => ATT1_n_308);
  ATT1_g13860 : NR2XD0BWP7T port map(A1 => ATT1_n_295, A2 => ATT1_n_285, ZN => ATT1_n_307);
  ATT1_g13861 : OAI21D0BWP7T port map(A1 => ATT1_n_285, A2 => ATT1_n_249, B => ATT1_n_302, ZN => ATT1_n_305);
  ATT1_g13862 : AOI21D0BWP7T port map(A1 => ATT1_n_298, A2 => ATT1_n_95, B => ATT1_n_97, ZN => ATT1_n_304);
  ATT1_g13863 : MAOI22D0BWP7T port map(A1 => ATT1_n_297, A2 => ATT1_n_106, B1 => ATT1_n_297, B2 => ATT1_n_106, ZN => ATT1_n_303);
  ATT1_g13864 : INVD0BWP7T port map(I => ATT1_n_295, ZN => ATT1_n_302);
  ATT1_g13865 : ND3D0BWP7T port map(A1 => ATT1_n_293, A2 => ATT1_n_271, A3 => ATT1_n_227, ZN => char1perctemp(4));
  ATT1_g13866 : INVD1BWP7T port map(I => FE_OFN2_ATT1_n_301, ZN => ATT1_n_300);
  ATT1_g13867 : OAI211D1BWP7T port map(A1 => ATT1_n_110, A2 => ATT1_n_287, B => ATT1_n_284, C => ATT1_n_137, ZN => ATT1_n_299);
  ATT1_g13868 : INR4D0BWP7T port map(A1 => ATT1_n_288, B1 => ATT1_n_118, B2 => ATT1_n_161, B3 => ATT1_n_284, ZN => ATT1_n_301);
  ATT1_g13869 : AO221D0BWP7T port map(A1 => ATT1_n_276, A2 => ATT1_n_191, B1 => ATT1_PM3_state1_0, B2 => char1perc(6), C => ATT1_n_202, Z => char1perctemp(6));
  ATT1_g13870 : OAI222D0BWP7T port map(A1 => ATT1_n_283, A2 => FE_DBTN13_char1perc_5, B1 => char1perc(5), B2 => ATT1_n_280, C1 => ATT1_n_199, C2 => ATT1_n_187, ZN => char1perctemp(5));
  ATT1_g13871 : OAI21D0BWP7T port map(A1 => ATT1_n_286, A2 => ATT1_n_77, B => ATT1_n_78, ZN => ATT1_n_298);
  ATT1_g13872 : AOI22D0BWP7T port map(A1 => ATT1_n_287, A2 => ATT1_n_137, B1 => ATT1_n_114, B2 => ATT1_n_129, ZN => ATT1_n_294);
  ATT1_g13873 : MOAI22D0BWP7T port map(A1 => ATT1_n_292, A2 => char2posy(5), B1 => ATT1_n_292, B2 => char2posy(5), ZN => ATT1_n_297);
  ATT1_g13874 : MAOI22D0BWP7T port map(A1 => ATT1_n_290, A2 => ATT1_n_107, B1 => ATT1_n_290, B2 => ATT1_n_107, ZN => ATT1_n_296);
  ATT1_g13875 : MAOI222D1BWP7T port map(A => ATT1_n_290, B => ATT1_n_68, C => char1posx(8), ZN => ATT1_n_295);
  ATT1_g13876 : ND3D0BWP7T port map(A1 => ATT1_n_277, A2 => ATT1_n_253, A3 => ATT1_n_228, ZN => char2perctemp(4));
  ATT1_g13877 : OAI221D0BWP7T port map(A1 => ATT1_n_269, A2 => ATT1_n_206, B1 => ATT1_n_101, B2 => ATT1_n_201, C => ATT1_n_209, ZN => char1perctemp(3));
  ATT1_g13878 : AOI21D0BWP7T port map(A1 => ATT1_n_281, A2 => char1perc(4), B => ATT1_n_219, ZN => ATT1_n_293);
  ATT1_g13879 : OAI211D1BWP7T port map(A1 => char1posy(4), A2 => ATT1_n_235, B => ATT1_n_251, C => ATT1_n_96, ZN => ATT1_n_292);
  ATT1_g13880 : OA221D0BWP7T port map(A1 => ATT1_n_237, A2 => ATT1_n_214, B1 => ATT1_n_135, B2 => ATT1_n_230, C => ATT1_n_279, Z => ATT1_n_291);
  ATT1_g13881 : AOI21D0BWP7T port map(A1 => ATT1_n_272, A2 => char2posx(7), B => ATT1_n_273, ZN => ATT1_n_290);
  ATT1_g13882 : NR2D1BWP7T port map(A1 => ATT1_n_278, A2 => ATT1_n_232, ZN => ATT1_n_289);
  ATT1_g13883 : NR2XD0BWP7T port map(A1 => ATT1_n_278, A2 => ATT1_n_233, ZN => ATT1_n_288);
  ATT1_g13884 : CKND1BWP7T port map(I => ATT1_n_287, ZN => ATT1_n_286);
  ATT1_g13885 : OA211D0BWP7T port map(A1 => FE_DBTN12_char1perc_4, A2 => ATT1_n_206, B => ATT1_n_275, C => ATT1_n_227, Z => ATT1_n_283);
  ATT1_g13886 : OAI222D0BWP7T port map(A1 => ATT1_n_274, A2 => FE_DBTN9_char2perc_5, B1 => char2perc(5), B2 => ATT1_n_259, C1 => ATT1_n_164, C2 => ATT1_n_189, ZN => char2perctemp(5));
  ATT1_g13887 : AOI21D0BWP7T port map(A1 => ATT1_n_233, A2 => ATT1_n_161, B => ATT1_n_278, ZN => ATT1_n_282);
  ATT1_g13888 : MAOI222D1BWP7T port map(A => ATT1_n_256, B => ATT1_n_53, C => char1posy(5), ZN => ATT1_n_287);
  ATT1_g13889 : OR4D1BWP7T port map(A1 => ATT1_n_162, A2 => ATT1_n_197, A3 => ATT1_n_237, A4 => ATT1_n_279, Z => ATT1_n_285);
  ATT1_g13890 : MOAI22D0BWP7T port map(A1 => ATT1_n_262, A2 => char2posy(4), B1 => ATT1_n_262, B2 => char2posy(4), ZN => ATT1_n_284);
  ATT1_g13891 : OAI221D0BWP7T port map(A1 => ATT1_n_247, A2 => ATT1_n_205, B1 => ATT1_n_102, B2 => ATT1_n_203, C => ATT1_n_211, ZN => char2perctemp(3));
  ATT1_g13892 : OAI221D0BWP7T port map(A1 => ATT1_n_201, A2 => ATT1_n_91, B1 => ATT1_n_139, B2 => ATT1_n_187, C => ATT1_n_275, ZN => ATT1_n_281);
  ATT1_g13893 : AO221D0BWP7T port map(A1 => ATT1_n_245, A2 => ATT1_n_190, B1 => ATT1_PM3_state2_0, B2 => char2perc(6), C => ATT1_n_204, Z => char2perctemp(6));
  ATT1_g13894 : OAI221D0BWP7T port map(A1 => ATT1_n_246, A2 => ATT1_n_206, B1 => char1perc(2), B2 => ATT1_n_201, C => ATT1_n_208, ZN => char1perctemp(2));
  ATT1_g13895 : OA21D0BWP7T port map(A1 => ATT1_n_201, A2 => ATT1_n_142, B => ATT1_n_271, Z => ATT1_n_280);
  ATT1_g13896 : MOAI22D0BWP7T port map(A1 => ATT1_n_260, A2 => char1perc(1), B1 => ATT1_n_265, B2 => char1perc(1), ZN => char1perctemp(1));
  ATT1_g13897 : AOI21D0BWP7T port map(A1 => ATT1_n_263, A2 => char2perc(4), B => ATT1_n_220, ZN => ATT1_n_277);
  ATT1_g13898 : MOAI22D0BWP7T port map(A1 => ATT1_n_268, A2 => char1perc(6), B1 => ATT1_n_268, B2 => char1perc(6), ZN => ATT1_n_276);
  ATT1_g13899 : MAOI22D0BWP7T port map(A1 => ATT1_n_261, A2 => ATT1_n_109, B1 => ATT1_n_261, B2 => ATT1_n_109, ZN => ATT1_n_279);
  ATT1_g13900 : XOR4D1BWP7T port map(A1 => ATT1_n_238, A2 => char2posy(2), A3 => char2posy(3), A4 => char1posy(3), Z => ATT1_n_278);
  ATT1_g13901 : OA211D0BWP7T port map(A1 => FE_DBTN8_char2perc_4, A2 => ATT1_n_205, B => ATT1_n_254, C => ATT1_n_228, Z => ATT1_n_274);
  ATT1_g13902 : AOI21D0BWP7T port map(A1 => ATT1_n_255, A2 => ATT1_n_89, B => char1posx(7), ZN => ATT1_n_273);
  ATT1_g13903 : ND3D0BWP7T port map(A1 => ATT1_n_255, A2 => ATT1_n_89, A3 => char1posx(7), ZN => ATT1_n_272);
  ATT1_g13904 : IAO21D0BWP7T port map(A1 => ATT1_n_252, A2 => ATT1_n_206, B => ATT1_PM3_state1_0, ZN => ATT1_n_275);
  ATT1_g13905 : AO32D1BWP7T port map(A1 => ATT1_n_242, A2 => ATT1_n_169, A3 => ATT1_PM3_state1_1, B1 => ATT1_PM3_state1_0, B2 => char1perc(7), Z => char1perctemp(7));
  ATT1_g13906 : OA21D0BWP7T port map(A1 => ATT1_n_248, A2 => ATT1_n_121, B => ATT1_n_266, Z => ATT1_n_270);
  ATT1_g13907 : MAOI22D0BWP7T port map(A1 => ATT1_n_244, A2 => ATT1_n_242, B1 => ATT1_n_242, B2 => char1perc(3), ZN => ATT1_n_269);
  ATT1_g13908 : IND3D1BWP7T port map(A1 => ATT1_n_206, B1 => FE_DBTN12_char1perc_4, B2 => ATT1_n_252, ZN => ATT1_n_271);
  ATT1_g13909 : AO211D0BWP7T port map(A1 => ATT1_n_191, A2 => ATT1_n_225, B => ATT1_n_202, C => ATT1_PM3_state1_0, Z => ATT1_n_265);
  ATT1_g13910 : OAI221D0BWP7T port map(A1 => ATT1_n_205, A2 => ATT1_n_213, B1 => char2perc(2), B2 => ATT1_n_203, C => ATT1_n_215, ZN => char2perctemp(2));
  ATT1_g13911 : NR2D0BWP7T port map(A1 => ATT1_n_249, A2 => ATT1_n_195, ZN => ATT1_n_264);
  ATT1_g13912 : OAI221D0BWP7T port map(A1 => ATT1_n_203, A2 => ATT1_n_75, B1 => ATT1_n_131, B2 => ATT1_n_189, C => ATT1_n_254, ZN => ATT1_n_263);
  ATT1_g13913 : OA221D0BWP7T port map(A1 => ATT1_n_226, A2 => ATT1_n_120, B1 => ATT1_n_79, B2 => ATT1_n_225, C => ATT1_n_243, Z => ATT1_n_268);
  ATT1_g13914 : ND2D1BWP7T port map(A1 => ATT1_n_249, A2 => ATT1_n_178, ZN => ATT1_n_267);
  ATT1_g13915 : ND2D1BWP7T port map(A1 => ATT1_n_249, A2 => ATT1_n_179, ZN => ATT1_n_266);
  ATT1_g13916 : AOI31D0BWP7T port map(A1 => ATT1_n_226, A2 => ATT1_n_169, A3 => ATT1_PM3_state1_1, B => ATT1_n_186, ZN => ATT1_n_260);
  ATT1_g13917 : MOAI22D0BWP7T port map(A1 => ATT1_n_231, A2 => char2perc(1), B1 => ATT1_n_240, B2 => char2perc(1), ZN => char2perctemp(1));
  ATT1_g13918 : OA21D0BWP7T port map(A1 => ATT1_n_203, A2 => ATT1_n_143, B => ATT1_n_253, Z => ATT1_n_259);
  ATT1_g13919 : MAOI22D0BWP7T port map(A1 => ATT1_n_241, A2 => ATT1_n_134, B1 => ATT1_n_241, B2 => ATT1_n_135, ZN => ATT1_n_258);
  ATT1_g13920 : MAOI22D0BWP7T port map(A1 => ATT1_n_241, A2 => ATT1_n_135, B1 => ATT1_n_241, B2 => ATT1_n_130, ZN => ATT1_n_257);
  ATT1_g13921 : MAOI22D0BWP7T port map(A1 => ATT1_n_235, A2 => ATT1_n_66, B1 => ATT1_n_235, B2 => ATT1_n_66, ZN => ATT1_n_262);
  ATT1_g13922 : MOAI22D0BWP7T port map(A1 => ATT1_n_236, A2 => char2posx(5), B1 => ATT1_n_236, B2 => char2posx(5), ZN => ATT1_n_261);
  ATT1_g13923 : AOI22D0BWP7T port map(A1 => ATT1_n_234, A2 => ATT1_n_96, B1 => ATT1_n_66, B2 => char2posy(4), ZN => ATT1_n_256);
  ATT1_g13924 : ND2D1BWP7T port map(A1 => ATT1_n_235, A2 => char2posy(4), ZN => ATT1_n_251);
  ATT1_g13925 : IOA21D1BWP7T port map(A1 => ATT1_n_161, A2 => ATT1_n_118, B => ATT1_n_232, ZN => ATT1_n_250);
  ATT1_g13926 : OR2D1BWP7T port map(A1 => ATT1_n_241, A2 => ATT1_n_90, Z => ATT1_n_255);
  ATT1_g13927 : IAO21D0BWP7T port map(A1 => ATT1_n_229, A2 => ATT1_n_205, B => ATT1_PM3_state2_0, ZN => ATT1_n_254);
  ATT1_g13928 : IND3D1BWP7T port map(A1 => ATT1_n_205, B1 => FE_DBTN8_char2perc_4, B2 => ATT1_n_229, ZN => ATT1_n_253);
  ATT1_g13929 : INR2D1BWP7T port map(A1 => ATT1_n_243, B1 => ATT1_n_239, ZN => ATT1_n_252);
  ATT1_g13930 : INVD1BWP7T port map(I => ATT1_n_249, ZN => ATT1_n_248);
  ATT1_g13931 : AO32D1BWP7T port map(A1 => ATT1_n_207, A2 => ATT1_n_168, A3 => ATT1_PM3_state2_1, B1 => ATT1_PM3_state2_0, B2 => char2perc(7), Z => char2perctemp(7));
  ATT1_g13932 : MAOI22D0BWP7T port map(A1 => ATT1_n_212, A2 => ATT1_n_207, B1 => ATT1_n_207, B2 => char2perc(3), ZN => ATT1_n_247);
  ATT1_g13933 : AOI22D0BWP7T port map(A1 => ATT1_n_226, A2 => ATT1_n_104, B1 => ATT1_n_225, B2 => char1perc(2), ZN => ATT1_n_246);
  ATT1_g13934 : MOAI22D0BWP7T port map(A1 => ATT1_n_216, A2 => char2perc(6), B1 => ATT1_n_216, B2 => char2perc(6), ZN => ATT1_n_245);
  ATT1_g13935 : OAI22D0BWP7T port map(A1 => ATT1_n_225, A2 => ATT1_n_150, B1 => ATT1_n_226, B2 => FE_DBTN11_char1perc_3, ZN => ATT1_n_244);
  ATT1_g13936 : MAOI22D0BWP7T port map(A1 => ATT1_n_217, A2 => ATT1_n_108, B1 => ATT1_n_217, B2 => ATT1_n_108, ZN => ATT1_n_249);
  ATT1_g13937 : OAI31D0BWP7T port map(A1 => char1perc(6), A2 => ATT1_n_74, A3 => ATT1_n_182, B => ATT1_n_222, ZN => char1percin(6));
  ATT1_g13938 : AO211D0BWP7T port map(A1 => ATT1_n_190, A2 => ATT1_n_184, B => ATT1_n_204, C => ATT1_PM3_state2_0, Z => ATT1_n_240);
  ATT1_g13939 : OAI31D0BWP7T port map(A1 => char2perc(7), A2 => ATT1_n_115, A3 => ATT1_n_163, B => ATT1_n_218, ZN => char2percin(7));
  ATT1_g13940 : OAI31D0BWP7T port map(A1 => char2perc(6), A2 => ATT1_n_92, A3 => ATT1_n_163, B => ATT1_n_223, ZN => char2percin(6));
  ATT1_g13941 : AOI21D0BWP7T port map(A1 => ATT1_n_128, A2 => FE_DBTN11_char1perc_3, B => ATT1_n_226, ZN => ATT1_n_239);
  ATT1_g13942 : OAI31D0BWP7T port map(A1 => char1perc(7), A2 => ATT1_n_116, A3 => ATT1_n_182, B => ATT1_n_221, ZN => char1percin(7));
  ATT1_g13943 : IND3D1BWP7T port map(A1 => ATT1_n_91, B1 => char1perc(1), B2 => ATT1_n_226, ZN => ATT1_n_243);
  ATT1_g13944 : OAI211D1BWP7T port map(A1 => char1posy(2), A2 => ATT1_n_160, B => ATT1_n_172, C => ATT1_n_80, ZN => ATT1_n_238);
  ATT1_g13945 : ND2D1BWP7T port map(A1 => ATT1_n_225, A2 => ATT1_n_128, ZN => ATT1_n_242);
  ATT1_g13946 : NR2XD0BWP7T port map(A1 => ATT1_n_210, A2 => ATT1_n_73, ZN => ATT1_n_241);
  ATT1_g13947 : INVD0BWP7T port map(I => ATT1_n_235, ZN => ATT1_n_234);
  ATT1_g13948 : INVD1BWP7T port map(I => ATT1_n_233, ZN => ATT1_n_232);
  ATT1_g13949 : AOI31D0BWP7T port map(A1 => ATT1_n_185, A2 => ATT1_n_168, A3 => ATT1_PM3_state2_1, B => ATT1_n_188, ZN => ATT1_n_231);
  ATT1_g13950 : INR3D0BWP7T port map(A1 => ATT1_n_197, B1 => ATT1_n_73, B2 => ATT1_n_134, ZN => ATT1_n_230);
  ATT1_g13951 : OAI222D0BWP7T port map(A1 => ATT1_n_176, A2 => ATT1_n_43, B1 => ATT1_n_62, B2 => ATT1_n_199, C1 => FE_DBTN13_char1perc_5, C2 => ATT1_n_166, ZN => char1percin(5));
  ATT1_g13952 : AO222D0BWP7T port map(A1 => ATT1_n_177, A2 => ATT1_PM3_state1_0, B1 => ATT1_n_150, B2 => ATT1_PM3_state1_1, C1 => ATT1_n_87, C2 => char1perc(3), Z => char1percin(3));
  ATT1_g13953 : OAI222D0BWP7T port map(A1 => ATT1_n_174, A2 => ATT1_n_44, B1 => ATT1_n_47, B2 => ATT1_n_157, C1 => FE_DBTN7_char2perc_3, C2 => ATT1_n_818, ZN => char2percin(3));
  ATT1_g13954 : OAI222D0BWP7T port map(A1 => ATT1_n_175, A2 => ATT1_n_44, B1 => ATT1_n_47, B2 => ATT1_n_164, C1 => FE_DBTN9_char2perc_5, C2 => ATT1_n_167, ZN => char2percin(5));
  ATT1_g13955 : OAI22D0BWP7T port map(A1 => ATT1_n_181, A2 => ATT1_n_111, B1 => ATT1_n_200, B2 => char1posx(4), ZN => ATT1_n_237);
  ATT1_g13956 : AOI31D0BWP7T port map(A1 => ATT1_n_180, A2 => char2posx(4), A3 => char1posx(4), B => ATT1_n_224, ZN => ATT1_n_236);
  ATT1_g13957 : MAOI222D1BWP7T port map(A => ATT1_n_173, B => FE_DBTN2_char1posy_3, C => char2posy(3), ZN => ATT1_n_235);
  ATT1_g13958 : MOAI22D0BWP7T port map(A1 => ATT1_n_183, A2 => char1posy(2), B1 => ATT1_n_183, B2 => char1posy(2), ZN => ATT1_n_233);
  ATT1_g13959 : INVD1BWP7T port map(I => ATT1_n_226, ZN => ATT1_n_225);
  ATT1_g13960 : NR3D0BWP7T port map(A1 => ATT1_n_180, A2 => char1posx(4), A3 => char2posx(4), ZN => ATT1_n_224);
  ATT1_g13961 : OAI21D0BWP7T port map(A1 => ATT1_n_193, A2 => ATT1_n_92, B => char2perc(6), ZN => ATT1_n_223);
  ATT1_g13962 : OAI21D0BWP7T port map(A1 => ATT1_n_192, A2 => ATT1_n_74, B => char1perc(6), ZN => ATT1_n_222);
  ATT1_g13963 : OAI21D0BWP7T port map(A1 => ATT1_n_192, A2 => ATT1_n_116, B => char1perc(7), ZN => ATT1_n_221);
  ATT1_g13964 : NR3D0BWP7T port map(A1 => ATT1_n_189, A2 => ATT1_n_132, A3 => char2perc(4), ZN => ATT1_n_220);
  ATT1_g13965 : AN3D0BWP7T port map(A1 => ATT1_n_186, A2 => ATT1_n_139, A3 => FE_DBTN12_char1perc_4, Z => ATT1_n_219);
  ATT1_g13966 : OAI21D0BWP7T port map(A1 => ATT1_n_193, A2 => ATT1_n_115, B => char2perc(7), ZN => ATT1_n_218);
  ATT1_g13967 : AOI21D0BWP7T port map(A1 => ATT1_n_184, A2 => ATT1_n_138, B => ATT1_n_140, ZN => ATT1_n_229);
  ATT1_g13968 : ND2D1BWP7T port map(A1 => ATT1_n_204, A2 => ATT1_n_143, ZN => ATT1_n_228);
  ATT1_g13969 : ND2D1BWP7T port map(A1 => ATT1_n_202, A2 => ATT1_n_142, ZN => ATT1_n_227);
  ATT1_g13970 : OAI31D1BWP7T port map(A1 => char1perc(6), A2 => char1perc(5), A3 => ATT1_n_170, B => char1perc(7), ZN => ATT1_n_226);
  ATT1_g13971 : AOI22D0BWP7T port map(A1 => ATT1_n_188, A2 => ATT1_n_105, B1 => char2perc(2), B2 => ATT1_PM3_state2_0, ZN => ATT1_n_215);
  ATT1_g13972 : OA21D0BWP7T port map(A1 => ATT1_n_133, A2 => ATT1_n_73, B => ATT1_n_197, Z => ATT1_n_214);
  ATT1_g13973 : MOAI22D0BWP7T port map(A1 => ATT1_n_182, A2 => char1perc(4), B1 => ATT1_n_192, B2 => char1perc(4), ZN => char1percin(4));
  ATT1_g13974 : AOI22D0BWP7T port map(A1 => ATT1_n_185, A2 => ATT1_n_105, B1 => ATT1_n_184, B2 => char2perc(2), ZN => ATT1_n_213);
  ATT1_g13975 : MOAI22D0BWP7T port map(A1 => ATT1_n_185, A2 => FE_DBTN7_char2perc_3, B1 => ATT1_n_185, B2 => ATT1_n_157, ZN => ATT1_n_212);
  ATT1_g13976 : MAOI22D0BWP7T port map(A1 => char2perc(3), A2 => ATT1_PM3_state2_0, B1 => ATT1_n_189, B2 => ATT1_n_157, ZN => ATT1_n_211);
  ATT1_g13977 : OAI31D0BWP7T port map(A1 => ATT1_n_82, A2 => ATT1_n_99, A3 => ATT1_n_181, B => ATT1_n_123, ZN => ATT1_n_210);
  ATT1_g13978 : AOI22D0BWP7T port map(A1 => ATT1_n_186, A2 => ATT1_n_150, B1 => char1perc(3), B2 => ATT1_PM3_state1_0, ZN => ATT1_n_209);
  ATT1_g13979 : AOI22D0BWP7T port map(A1 => ATT1_n_186, A2 => ATT1_n_104, B1 => char1perc(2), B2 => ATT1_PM3_state1_0, ZN => ATT1_n_208);
  ATT1_g13980 : MOAI22D0BWP7T port map(A1 => ATT1_n_163, A2 => char2perc(4), B1 => ATT1_n_193, B2 => char2perc(4), ZN => char2percin(4));
  ATT1_g13981 : MOAI22D0BWP7T port map(A1 => ATT1_n_194, A2 => char2posx(3), B1 => ATT1_n_194, B2 => char2posx(3), ZN => ATT1_n_217);
  ATT1_g13982 : AOI22D0BWP7T port map(A1 => ATT1_n_185, A2 => ATT1_n_152, B1 => ATT1_n_184, B2 => ATT1_n_119, ZN => ATT1_n_216);
  ATT1_g13983 : INVD0BWP7T port map(I => ATT1_n_204, ZN => ATT1_n_203);
  ATT1_g13984 : INVD1BWP7T port map(I => ATT1_n_202, ZN => ATT1_n_201);
  ATT1_g13985 : ND2D1BWP7T port map(A1 => ATT1_n_181, A2 => char2posx(4), ZN => ATT1_n_200);
  ATT1_g13986 : ND2D1BWP7T port map(A1 => ATT1_n_184, A2 => ATT1_n_127, ZN => ATT1_n_207);
  ATT1_g13987 : ND2D1BWP7T port map(A1 => ATT1_n_191, A2 => ATT1_n_169, ZN => ATT1_n_206);
  ATT1_g13988 : ND2D1BWP7T port map(A1 => ATT1_n_190, A2 => ATT1_n_168, ZN => ATT1_n_205);
  ATT1_g13989 : INR2XD0BWP7T port map(A1 => ATT1_n_190, B1 => ATT1_n_168, ZN => ATT1_n_204);
  ATT1_g13990 : INR2XD0BWP7T port map(A1 => ATT1_n_191, B1 => ATT1_n_169, ZN => ATT1_n_202);
  ATT1_g13991 : INVD0BWP7T port map(I => ATT1_n_195, ZN => ATT1_n_196);
  ATT1_g13992 : AO222D0BWP7T port map(A1 => ATT1_n_146, A2 => ATT1_PM3_state2_0, B1 => ATT1_n_105, B2 => ATT1_PM3_state2_1, C1 => ATT1_n_71, C2 => char2perc(2), Z => char2percin(2));
  ATT1_g13993 : AO222D0BWP7T port map(A1 => ATT1_n_147, A2 => ATT1_PM3_state1_0, B1 => ATT1_n_104, B2 => ATT1_PM3_state1_1, C1 => ATT1_n_87, C2 => char1perc(2), Z => char1percin(2));
  ATT1_g13994 : MAOI22D0BWP7T port map(A1 => ATT1_n_170, A2 => FE_DBTN13_char1perc_5, B1 => ATT1_n_170, B2 => FE_DBTN13_char1perc_5, ZN => ATT1_n_199);
  ATT1_g13995 : INR2D1BWP7T port map(A1 => ATT1_n_121, B1 => ATT1_n_179, ZN => ATT1_n_198);
  ATT1_g13996 : INR2XD0BWP7T port map(A1 => ATT1_n_82, B1 => ATT1_n_180, ZN => ATT1_n_197);
  ATT1_g13997 : NR2XD0BWP7T port map(A1 => ATT1_n_178, A2 => ATT1_n_121, ZN => ATT1_n_195);
  ATT1_g13998 : CKND1BWP7T port map(I => ATT1_n_189, ZN => ATT1_n_188);
  ATT1_g13999 : INVD0BWP7T port map(I => ATT1_n_187, ZN => ATT1_n_186);
  ATT1_g14000 : INVD1BWP7T port map(I => ATT1_n_185, ZN => ATT1_n_184);
  ATT1_g14001 : AOI211XD0BWP7T port map(A1 => ATT1_n_124, A2 => char2posx(2), B => ATT1_n_158, C => ATT1_n_85, ZN => ATT1_n_194);
  ATT1_g14002 : ND2D1BWP7T port map(A1 => ATT1_n_167, A2 => ATT1_n_131, ZN => ATT1_n_193);
  ATT1_g14003 : ND2D1BWP7T port map(A1 => ATT1_n_166, A2 => ATT1_n_139, ZN => ATT1_n_192);
  ATT1_g14004 : NR2XD0BWP7T port map(A1 => ATT1_n_165, A2 => ATT1_n_62, ZN => ATT1_n_191);
  ATT1_g14005 : NR2XD0BWP7T port map(A1 => ATT1_n_171, A2 => ATT1_n_47, ZN => ATT1_n_190);
  ATT1_g14006 : ND2D1BWP7T port map(A1 => ATT1_n_171, A2 => ATT1_PM3_state2_1, ZN => ATT1_n_189);
  ATT1_g14007 : ND2D1BWP7T port map(A1 => ATT1_n_165, A2 => ATT1_PM3_state1_1, ZN => ATT1_n_187);
  ATT1_g14008 : OAI31D0BWP7T port map(A1 => char2perc(6), A2 => char2perc(5), A3 => ATT1_n_154, B => char2perc(7), ZN => ATT1_n_185);
  ATT1_g14009 : INVD0BWP7T port map(I => ATT1_n_181, ZN => ATT1_n_180);
  ATT1_g14010 : INVD1BWP7T port map(I => ATT1_n_179, ZN => ATT1_n_178);
  ATT1_g14011 : MOAI22D0BWP7T port map(A1 => ATT1_n_141, A2 => FE_DBTN11_char1perc_3, B1 => ATT1_n_141, B2 => FE_DBTN11_char1perc_3, ZN => ATT1_n_177);
  ATT1_g14012 : AOI32D1BWP7T port map(A1 => ATT1_n_155, A2 => FE_DBTN13_char1perc_5, A3 => char1perc(4), B1 => FE_DBTN12_char1perc_4, B2 => char1perc(5), ZN => ATT1_n_176);
  ATT1_g14013 : AOI32D1BWP7T port map(A1 => ATT1_n_156, A2 => FE_DBTN9_char2perc_5, A3 => char2perc(4), B1 => FE_DBTN8_char2perc_4, B2 => char2perc(5), ZN => ATT1_n_175);
  ATT1_g14014 : MAOI22D0BWP7T port map(A1 => ATT1_n_136, A2 => FE_DBTN7_char2perc_3, B1 => ATT1_n_136, B2 => FE_DBTN7_char2perc_3, ZN => ATT1_n_174);
  ATT1_g14015 : MOAI22D0BWP7T port map(A1 => ATT1_n_49, A2 => char1posy(2), B1 => ATT1_n_160, B2 => ATT1_n_80, ZN => ATT1_n_173);
  ATT1_g14016 : OA21D0BWP7T port map(A1 => ATT1_n_160, A2 => char2posy(2), B => ATT1_n_172, Z => ATT1_n_183);
  ATT1_g14017 : AOI22D0BWP7T port map(A1 => ATT1_n_155, A2 => ATT1_PM3_state1_0, B1 => ATT1_n_139, B2 => ATT1_PM3_state1_1, ZN => ATT1_n_182);
  ATT1_g14018 : MAOI222D1BWP7T port map(A => ATT1_n_144, B => ATT1_n_67, C => char2posx(3), ZN => ATT1_n_181);
  ATT1_g14019 : MAOI22D0BWP7T port map(A1 => ATT1_n_159, A2 => char2posx(2), B1 => ATT1_n_159, B2 => char2posx(2), ZN => ATT1_n_179);
  ATT1_g14020 : ND2D1BWP7T port map(A1 => ATT1_n_160, A2 => char2posy(2), ZN => ATT1_n_172);
  ATT1_g14021 : NR3D0BWP7T port map(A1 => ATT1_n_153, A2 => char2perc(6), A3 => char2perc(7), ZN => ATT1_n_171);
  ATT1_g14022 : AN2D0BWP7T port map(A1 => ATT1_n_139, A2 => char1perc(4), Z => ATT1_n_170);
  ATT1_g14023 : IND3D1BWP7T port map(A1 => char1perc(7), B1 => ATT1_n_116, B2 => ATT1_n_145, ZN => ATT1_n_169);
  ATT1_g14024 : IND3D1BWP7T port map(A1 => char2perc(7), B1 => ATT1_n_115, B2 => ATT1_n_148, ZN => ATT1_n_168);
  ATT1_g14025 : AO211D0BWP7T port map(A1 => ATT1_n_122, A2 => ATT1_n_123, B => ATT1_n_149, C => ATT1_n_126, Z => ATT1_n_162);
  ATT1_g14026 : OA21D0BWP7T port map(A1 => ATT1_n_156, A2 => ATT1_n_44, B => ATT1_n_818, Z => ATT1_n_167);
  ATT1_g14027 : OA21D0BWP7T port map(A1 => ATT1_n_155, A2 => ATT1_n_43, B => ATT1_n_828, Z => ATT1_n_166);
  ATT1_g14028 : NR3D0BWP7T port map(A1 => ATT1_n_151, A2 => char1perc(6), A3 => char1perc(7), ZN => ATT1_n_165);
  ATT1_g14029 : MAOI22D0BWP7T port map(A1 => ATT1_n_154, A2 => FE_DBTN9_char2perc_5, B1 => ATT1_n_154, B2 => FE_DBTN9_char2perc_5, ZN => ATT1_n_164);
  ATT1_g14030 : AOI22D0BWP7T port map(A1 => ATT1_n_156, A2 => ATT1_PM3_state2_0, B1 => ATT1_n_131, B2 => ATT1_PM3_state2_1, ZN => ATT1_n_163);
  ATT1_g14031 : FA1D0BWP7T port map(A => ATT1_n_51, B => char2posy(1), CI => ATT1_n_86, CO => ATT1_n_160, S => ATT1_n_161);
  ATT1_g14032 : HA1D0BWP7T port map(A => ATT1_n_50, B => ATT1_n_125, CO => ATT1_n_158, S => ATT1_n_159);
  ATT1_g14033 : OAI222D0BWP7T port map(A1 => ATT1_n_103, A2 => ATT1_n_43, B1 => FE_DBTN10_char1perc_1, B2 => ATT1_n_828, C1 => ATT1_n_62, C2 => char1perc(1), ZN => char1percin(1));
  ATT1_g14034 : OAI222D0BWP7T port map(A1 => ATT1_n_100, A2 => ATT1_n_44, B1 => FE_DBTN5_char2perc_1, B2 => ATT1_n_818, C1 => char2perc(1), C2 => ATT1_n_47, ZN => char2percin(1));
  ATT1_g14035 : AOI21D0BWP7T port map(A1 => ATT1_n_84, A2 => FE_DBTN5_char2perc_1, B => ATT1_n_92, ZN => ATT1_n_153);
  ATT1_g14036 : IND2D1BWP7T port map(A1 => ATT1_n_140, B1 => ATT1_n_81, ZN => ATT1_n_152);
  ATT1_g14037 : AOI21D0BWP7T port map(A1 => ATT1_n_98, A2 => FE_DBTN10_char1perc_1, B => ATT1_n_74, ZN => ATT1_n_151);
  ATT1_g14038 : NR2XD0BWP7T port map(A1 => ATT1_n_140, A2 => ATT1_n_132, ZN => ATT1_n_157);
  ATT1_g14039 : OAI21D0BWP7T port map(A1 => ATT1_n_94, A2 => FE_DBTN7_char2perc_3, B => ATT1_n_75, ZN => ATT1_n_156);
  ATT1_g14040 : OAI21D0BWP7T port map(A1 => ATT1_n_93, A2 => FE_DBTN11_char1perc_3, B => ATT1_n_91, ZN => ATT1_n_155);
  ATT1_g14041 : NR2D1BWP7T port map(A1 => ATT1_n_132, A2 => FE_DBTN8_char2perc_4, ZN => ATT1_n_154);
  ATT1_g14042 : MOAI22D0BWP7T port map(A1 => ATT1_n_122, A2 => ATT1_n_72, B1 => ATT1_n_112, B2 => ATT1_n_89, ZN => ATT1_n_149);
  ATT1_g14043 : IND3D1BWP7T port map(A1 => ATT1_n_84, B1 => char2perc(5), B2 => char2perc(6), ZN => ATT1_n_148);
  ATT1_g14044 : OAI21D0BWP7T port map(A1 => ATT1_n_93, A2 => ATT1_n_58, B => ATT1_n_141, ZN => ATT1_n_147);
  ATT1_g14045 : OAI21D0BWP7T port map(A1 => ATT1_n_94, A2 => FE_DBTN6_char2perc_2, B => ATT1_n_136, ZN => ATT1_n_146);
  ATT1_g14046 : IND3D1BWP7T port map(A1 => ATT1_n_98, B1 => char1perc(5), B2 => char1perc(6), ZN => ATT1_n_145);
  ATT1_g14047 : MOAI22D0BWP7T port map(A1 => ATT1_n_125, A2 => ATT1_n_85, B1 => ATT1_n_50, B2 => char2posx(2), ZN => ATT1_n_144);
  ATT1_g14048 : MAOI22D0BWP7T port map(A1 => ATT1_n_76, A2 => char1perc(3), B1 => ATT1_n_76, B2 => char1perc(3), ZN => ATT1_n_150);
  ATT1_g14049 : ND2D1BWP7T port map(A1 => ATT1_n_127, A2 => FE_DBTN7_char2perc_3, ZN => ATT1_n_138);
  ATT1_g14050 : AN2D1BWP7T port map(A1 => ATT1_n_75, A2 => FE_DBTN8_char2perc_4, Z => ATT1_n_143);
  ATT1_g14051 : AN2D1BWP7T port map(A1 => ATT1_n_91, A2 => FE_DBTN12_char1perc_4, Z => ATT1_n_142);
  ATT1_g14052 : ND2D1BWP7T port map(A1 => ATT1_n_93, A2 => ATT1_n_58, ZN => ATT1_n_141);
  ATT1_g14053 : NR2D1BWP7T port map(A1 => ATT1_n_75, A2 => FE_DBTN5_char2perc_1, ZN => ATT1_n_140);
  ATT1_g14054 : ND2D1BWP7T port map(A1 => ATT1_n_76, A2 => FE_DBTN11_char1perc_3, ZN => ATT1_n_139);
  ATT1_g14055 : INVD1BWP7T port map(I => ATT1_n_134, ZN => ATT1_n_133);
  ATT1_g14056 : INVD1BWP7T port map(I => ATT1_n_132, ZN => ATT1_n_131);
  ATT1_g14057 : AOI22D0BWP7T port map(A1 => ATT1_n_112, A2 => ATT1_n_88, B1 => ATT1_n_113, B2 => ATT1_n_90, ZN => ATT1_n_130);
  ATT1_g14058 : IND2D1BWP7T port map(A1 => ATT1_n_114, B1 => ATT1_n_78, ZN => ATT1_n_137);
  ATT1_g14059 : ND2D1BWP7T port map(A1 => ATT1_n_94, A2 => FE_DBTN6_char2perc_2, ZN => ATT1_n_136);
  ATT1_g14060 : INR2XD0BWP7T port map(A1 => ATT1_n_89, B1 => ATT1_n_122, ZN => ATT1_n_135);
  ATT1_g14061 : AOI21D0BWP7T port map(A1 => ATT1_n_112, A2 => ATT1_n_90, B => ATT1_n_126, ZN => ATT1_n_134);
  ATT1_g14062 : AOI21D0BWP7T port map(A1 => char2perc(1), A2 => char2perc(2), B => char2perc(3), ZN => ATT1_n_132);
  ATT1_g14063 : INVD0BWP7T port map(I => ATT1_n_77, ZN => ATT1_n_129);
  ATT1_g14064 : INVD0BWP7T port map(I => ATT1_n_125, ZN => ATT1_n_124);
  ATT1_g14065 : ND2D1BWP7T port map(A1 => ATT1_n_120, A2 => char1perc(6), ZN => ATT1_n_128);
  ATT1_g14066 : IND2D1BWP7T port map(A1 => ATT1_n_119, B1 => char2perc(6), ZN => ATT1_n_127);
  ATT1_g14067 : NR2D0BWP7T port map(A1 => ATT1_n_112, A2 => ATT1_n_89, ZN => ATT1_n_126);
  ATT1_g14068 : NR2D1BWP7T port map(A1 => ATT1_n_117, A2 => ATT1_n_83, ZN => ATT1_n_125);
  ATT1_g14069 : OAI222D0BWP7T port map(A1 => ATT1_PM3_state1_0, A2 => ATT1_n_65, B1 => ATT1_n_65, B2 => ATT1_n_62, C1 => char1perc(0), C2 => ATT1_n_43, ZN => char1percin(0));
  ATT1_g14070 : OAI222D0BWP7T port map(A1 => ATT1_PM3_state2_0, A2 => FE_DBTN4_char2perc_0, B1 => FE_DBTN4_char2perc_0, B2 => ATT1_n_47, C1 => char2perc(0), C2 => ATT1_n_44, ZN => char2percin(0));
  ATT1_g14071 : IND3D1BWP7T port map(A1 => ATT1_n_99, B1 => char2posx(4), B2 => FE_DBTN3_char1posx_4, ZN => ATT1_n_123);
  ATT1_g14072 : IND2D1BWP7T port map(A1 => ATT1_n_90, B1 => ATT1_n_113, ZN => ATT1_n_122);
  ATT1_g14073 : IND3D1BWP7T port map(A1 => ATT1_n_83, B1 => ATT1_n_70, B2 => ATT1_n_117, ZN => ATT1_n_121);
  ATT1_g14074 : INVD1BWP7T port map(I => ATT1_n_113, ZN => ATT1_n_112);
  ATT1_g14075 : NR2D0BWP7T port map(A1 => ATT1_n_87, A2 => ATT1_n_65, ZN => char1perctemp(0));
  ATT1_g14076 : MAOI22D0BWP7T port map(A1 => char2posx(4), A2 => char1posx(4), B1 => char2posx(4), B2 => char1posx(4), ZN => ATT1_n_111);
  ATT1_g14077 : NR2D0BWP7T port map(A1 => ATT1_n_71, A2 => FE_DBTN4_char2perc_0, ZN => char2perctemp(0));
  ATT1_g14078 : ND2D1BWP7T port map(A1 => ATT1_n_79, A2 => FE_DBTN11_char1perc_3, ZN => ATT1_n_120);
  ATT1_g14079 : CKAN2D1BWP7T port map(A1 => ATT1_n_81, A2 => FE_DBTN7_char2perc_3, Z => ATT1_n_119);
  ATT1_g14080 : MAOI22D0BWP7T port map(A1 => char2posy(0), A2 => char1posy(0), B1 => char2posy(0), B2 => char1posy(0), ZN => ATT1_n_118);
  ATT1_g14081 : AOI22D0BWP7T port map(A1 => FE_DBTN0_char2posx_0, A2 => char1posx(0), B1 => FE_DBTN1_char2posx_1, B2 => char1posx(1), ZN => ATT1_n_117);
  ATT1_g14082 : IND2D1BWP7T port map(A1 => ATT1_n_74, B1 => char1perc(6), ZN => ATT1_n_116);
  ATT1_g14083 : IND2D1BWP7T port map(A1 => ATT1_n_92, B1 => char2perc(6), ZN => ATT1_n_115);
  ATT1_g14084 : INR2XD0BWP7T port map(A1 => ATT1_n_95, B1 => ATT1_n_97, ZN => ATT1_n_114);
  ATT1_g14085 : MOAI22D0BWP7T port map(A1 => char1posx(7), A2 => char2posx(7), B1 => char2posx(7), B2 => char1posx(7), ZN => ATT1_n_113);
  ATT1_g14086 : AOI22D0BWP7T port map(A1 => char1perc(1), A2 => ATT1_n_65, B1 => FE_DBTN10_char1perc_1, B2 => char1perc(0), ZN => ATT1_n_103);
  ATT1_g14087 : AOI22D0BWP7T port map(A1 => FE_DBTN6_char2perc_2, A2 => char2perc(3), B1 => FE_DBTN7_char2perc_3, B2 => char2perc(2), ZN => ATT1_n_102);
  ATT1_g14088 : AOI22D0BWP7T port map(A1 => ATT1_n_58, A2 => char1perc(3), B1 => FE_DBTN11_char1perc_3, B2 => char1perc(2), ZN => ATT1_n_101);
  ATT1_g14089 : AOI22D0BWP7T port map(A1 => char2perc(1), A2 => FE_DBTN4_char2perc_0, B1 => FE_DBTN5_char2perc_1, B2 => char2perc(0), ZN => ATT1_n_100);
  ATT1_g14090 : MOAI22D0BWP7T port map(A1 => char1posy(6), A2 => char2posy(6), B1 => char2posy(6), B2 => char1posy(6), ZN => ATT1_n_110);
  ATT1_g14091 : MAOI22D0BWP7T port map(A1 => FE_DBTN3_char1posx_4, A2 => char1posx(5), B1 => FE_DBTN3_char1posx_4, B2 => char1posx(5), ZN => ATT1_n_109);
  ATT1_g14092 : MAOI22D0BWP7T port map(A1 => ATT1_n_67, A2 => char2posx(2), B1 => ATT1_n_67, B2 => char2posx(2), ZN => ATT1_n_108);
  ATT1_g14093 : MOAI22D0BWP7T port map(A1 => char1posx(8), A2 => FE_PHN123_char2posx_8, B1 => FE_PHN123_char2posx_8, B2 => char1posx(8), ZN => ATT1_n_107);
  ATT1_g14094 : MAOI22D0BWP7T port map(A1 => ATT1_n_66, A2 => char1posy(5), B1 => ATT1_n_66, B2 => char1posy(5), ZN => ATT1_n_106);
  ATT1_g14095 : OAI22D0BWP7T port map(A1 => FE_DBTN6_char2perc_2, A2 => char2perc(1), B1 => FE_DBTN5_char2perc_1, B2 => char2perc(2), ZN => ATT1_n_105);
  ATT1_g14096 : OAI22D0BWP7T port map(A1 => ATT1_n_58, A2 => char1perc(1), B1 => FE_DBTN10_char1perc_1, B2 => char1perc(2), ZN => ATT1_n_104);
  ATT1_g14097 : INVD0BWP7T port map(I => ATT1_n_89, ZN => ATT1_n_88);
  ATT1_g14098 : INVD0BWP7T port map(I => ATT1_n_87, ZN => ATT1_n_828);
  ATT1_g14099 : ND2D1BWP7T port map(A1 => ATT1_PM4_state2_1, A2 => ATT1_PM4_state2_0, ZN => char2death);
  ATT1_g14100 : INR2XD0BWP7T port map(A1 => char1posx(5), B1 => char2posx(5), ZN => ATT1_n_99);
  ATT1_g14101 : NR2XD0BWP7T port map(A1 => char1perc(2), A2 => char1perc(3), ZN => ATT1_n_98);
  ATT1_g14102 : INR2D1BWP7T port map(A1 => char2posy(7), B1 => char1posy(7), ZN => ATT1_n_97);
  ATT1_g14103 : AN2D1BWP7T port map(A1 => ATT1_PM2_state2_1, A2 => ATT1_PM2_state2_0, Z => ATT1_at2a);
  ATT1_g14104 : IND2D1BWP7T port map(A1 => char2posy(4), B1 => char1posy(4), ZN => ATT1_n_96);
  ATT1_g14105 : CKAN2D1BWP7T port map(A1 => FE_PHN116_ATT1_PM2_state1_1, A2 => ATT1_PM2_state1_0, Z => ATT1_at1a);
  ATT1_g14106 : IND2D1BWP7T port map(A1 => char2posy(7), B1 => char1posy(7), ZN => ATT1_n_95);
  ATT1_g14107 : ND2D1BWP7T port map(A1 => char2perc(1), A2 => char2perc(0), ZN => ATT1_n_94);
  ATT1_g14108 : IND2D1BWP7T port map(A1 => char2posy(0), B1 => char1posy(0), ZN => ATT1_n_86);
  ATT1_g14109 : ND2D1BWP7T port map(A1 => char1perc(1), A2 => char1perc(0), ZN => ATT1_n_93);
  ATT1_g14110 : ND2D1BWP7T port map(A1 => char2perc(4), A2 => char2perc(5), ZN => ATT1_n_92);
  ATT1_g14111 : CKND2D1BWP7T port map(A1 => char1perc(2), A2 => char1perc(3), ZN => ATT1_n_91);
  ATT1_g14112 : INR2XD0BWP7T port map(A1 => char1posx(6), B1 => char2posx(6), ZN => ATT1_n_90);
  ATT1_g14113 : IND2D1BWP7T port map(A1 => char1posx(6), B1 => char2posx(6), ZN => ATT1_n_89);
  ATT1_g14114 : NR2XD0BWP7T port map(A1 => ATT1_PM3_state1_1, A2 => ATT1_PM3_state1_0, ZN => ATT1_n_87);
  ATT1_g14115 : INVD0BWP7T port map(I => ATT1_n_73, ZN => ATT1_n_72);
  ATT1_g14116 : INVD1BWP7T port map(I => ATT1_n_71, ZN => ATT1_n_818);
  ATT1_g14117 : ND2D1BWP7T port map(A1 => ATT1_PM4_state1_1, A2 => ATT1_PM4_state1_0, ZN => char1death);
  ATT1_g14118 : IND2D1BWP7T port map(A1 => char1posx(0), B1 => char2posx(0), ZN => ATT1_n_70);
  ATT1_g14119 : NR2D1BWP7T port map(A1 => ATT1_n_50, A2 => char2posx(2), ZN => ATT1_n_85);
  ATT1_g14120 : NR2XD0BWP7T port map(A1 => char2perc(2), A2 => char2perc(3), ZN => ATT1_n_84);
  ATT1_g14121 : NR2XD0BWP7T port map(A1 => FE_DBTN1_char2posx_1, A2 => char1posx(1), ZN => ATT1_n_83);
  ATT1_g14122 : NR2XD0BWP7T port map(A1 => FE_DBTN3_char1posx_4, A2 => char2posx(4), ZN => ATT1_n_82);
  ATT1_g14123 : NR2XD0BWP7T port map(A1 => char2perc(5), A2 => char2perc(4), ZN => ATT1_n_81);
  ATT1_g14124 : ND2D1BWP7T port map(A1 => ATT1_n_49, A2 => char1posy(2), ZN => ATT1_n_80);
  ATT1_g14125 : NR2XD0BWP7T port map(A1 => char1perc(5), A2 => char1perc(4), ZN => ATT1_n_79);
  ATT1_g14126 : IND2D1BWP7T port map(A1 => char1posy(6), B1 => char2posy(6), ZN => ATT1_n_78);
  ATT1_g14127 : INR2D1BWP7T port map(A1 => char1posy(6), B1 => char2posy(6), ZN => ATT1_n_77);
  ATT1_g14128 : CKND2D1BWP7T port map(A1 => char1perc(2), A2 => char1perc(1), ZN => ATT1_n_76);
  ATT1_g14129 : CKND2D1BWP7T port map(A1 => char2perc(2), A2 => char2perc(3), ZN => ATT1_n_75);
  ATT1_g14130 : ND2D1BWP7T port map(A1 => char1perc(4), A2 => char1perc(5), ZN => ATT1_n_74);
  ATT1_g14131 : INR2D1BWP7T port map(A1 => char2posx(5), B1 => char1posx(5), ZN => ATT1_n_73);
  ATT1_g14132 : NR2XD0BWP7T port map(A1 => ATT1_PM3_state2_0, A2 => ATT1_PM3_state2_1, ZN => ATT1_n_71);
  ATT1_g14134 : INVD0BWP7T port map(I => FE_PHN123_char2posx_8, ZN => ATT1_n_68);
  ATT1_g14135 : INVD1BWP7T port map(I => char1posx(3), ZN => ATT1_n_67);
  ATT1_g14136 : INVD1BWP7T port map(I => char1posy(4), ZN => ATT1_n_66);
  ATT1_g14137 : INVD1BWP7T port map(I => char1perc(0), ZN => ATT1_n_65);
  ATT1_g14144 : INVD1BWP7T port map(I => char1perc(2), ZN => ATT1_n_58);
  ATT1_g14149 : INVD0BWP7T port map(I => char2posy(5), ZN => ATT1_n_53);
  ATT1_g14151 : CKND1BWP7T port map(I => char1posy(1), ZN => ATT1_n_51);
  ATT1_g14152 : INVD1BWP7T port map(I => char1posx(2), ZN => ATT1_n_50);
  ATT1_g14153 : CKND1BWP7T port map(I => char2posy(2), ZN => ATT1_n_49);
  ATT1_g2 : INR2D1BWP7T port map(A1 => ATT1_n_654, B1 => ATT1_n_598, ZN => ATT1_n_42);
  ATT1_g14160 : INR2D1BWP7T port map(A1 => ATT1_n_631, B1 => ATT1_n_705, ZN => ATT1_n_41);
  ATT1_g14161 : IND2D1BWP7T port map(A1 => ATT1_n_457, B1 => ATT1_n_336, ZN => ATT1_n_40);
  ATT1_g14162 : INR3D0BWP7T port map(A1 => ATT1_n_326, B1 => ATT1_n_317, B2 => ATT1_n_473, ZN => ATT1_n_39);
  ATT1_g14163 : INR3D0BWP7T port map(A1 => ATT1_n_319, B1 => ATT1_n_350, B2 => ATT1_n_323, ZN => ATT1_n_38);
  ATT1_PM4_state1_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => ATT1_n_36, Q => ATT1_PM4_state1_1);
  ATT1_PM4_state2_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_15, D => ATT1_n_37, Q => FE_PHN115_ATT1_PM4_state2_1);
  ATT1_PM2_state2_reg_1 : DFQD1BWP7T port map(CP => CTS_16, D => FE_PHN145_ATT1_n_35, Q => FE_PHN121_ATT1_PM2_state2_1);
  ATT1_PM2_state1_reg_1 : DFQD1BWP7T port map(CP => CTS_16, D => FE_PHN157_ATT1_n_34, Q => ATT1_PM2_state1_1);
  ATT1_PM2_state1_reg_0 : DFQD1BWP7T port map(CP => CTS_16, D => ATT1_n_32, Q => ATT1_PM2_state1_0);
  ATT1_PM2_state2_reg_0 : DFQD1BWP7T port map(CP => CTS_16, D => ATT1_n_33, Q => FE_PHN120_ATT1_PM2_state2_0);
  ATT1_g794 : OAI211D1BWP7T port map(A1 => char2posx(7), A2 => ATT1_n_28, B => ATT1_n_22, C => FE_PHN123_char2posx_8, ZN => ATT1_n_37);
  ATT1_g795 : OAI211D1BWP7T port map(A1 => char1posx(7), A2 => ATT1_n_29, B => ATT1_n_19, C => char1posx(8), ZN => ATT1_n_36);
  ATT1_g796 : AO221D0BWP7T port map(A1 => ATT1_n_11, A2 => FE_PHN98_inputsp2_5, B1 => ATT1_n_16, B2 => ATT1_PM2_state2_1, C => ATT1_n_31, Z => ATT1_n_35);
  ATT1_g797 : AO221D0BWP7T port map(A1 => ATT1_n_13, A2 => inputsp1(5), B1 => ATT1_at1a, B2 => ATT1_n_7, C => ATT1_n_30, Z => ATT1_n_34);
  ATT1_g798 : AO211D0BWP7T port map(A1 => ATT1_n_20, A2 => FE_DBTN14_reset, B => ATT1_n_0, C => ATT1_n_16, Z => ATT1_n_33);
  ATT1_g799 : AO22D0BWP7T port map(A1 => ATT1_n_27, A2 => FE_DBTN14_reset, B1 => ATT1_n_7, B2 => ATT1_PM2_state1_0, Z => FE_PHN148_ATT1_n_32);
  ATT1_PM2_state2_reg_2 : DFQD1BWP7T port map(CP => CTS_16, D => FE_PHN126_ATT1_n_25, Q => ATT1_at2b);
  ATT1_g802 : IAO21D0BWP7T port map(A1 => ATT1_n_21, A2 => ATT1_n_0, B => inputsp2(4), ZN => ATT1_n_31);
  ATT1_g803 : NR4D0BWP7T port map(A1 => ATT1_n_15, A2 => inputsp1(4), A3 => FE_PHN116_ATT1_PM2_state1_1, A4 => FE_OFN3_reset, ZN => ATT1_n_30);
  ATT1_g808 : INR3D0BWP7T port map(A1 => char1posx(4), B1 => ATT1_n_4, B2 => ATT1_n_8, ZN => ATT1_n_29);
  ATT1_g809 : INR3D0BWP7T port map(A1 => char2posx(4), B1 => ATT1_n_3, B2 => ATT1_n_9, ZN => ATT1_n_28);
  ATT1_g810 : IAO21D0BWP7T port map(A1 => ATT1_n_14, A2 => ATT1_PM2_state1_0, B => FE_PHN116_ATT1_PM2_state1_1, ZN => ATT1_n_27);
  ATT1_g811 : MOAI22D0BWP7T port map(A1 => FE_PHN146_ATT1_n_12, A2 => inputsp1(5), B1 => ATT1_at1b, B2 => ATT1_n_7, ZN => ATT1_n_26);
  ATT1_g812 : MOAI22D0BWP7T port map(A1 => ATT1_n_10, A2 => FE_PHN98_inputsp2_5, B1 => ATT1_at2b, B2 => ATT1_n_7, ZN => ATT1_n_25);
  ATT1_g813 : INR2XD0BWP7T port map(A1 => ATT1_n_18, B1 => ATT1_at2a, ZN => ATT1_n_24);
  ATT1_g814 : INR2XD0BWP7T port map(A1 => ATT1_n_17, B1 => ATT1_at1a, ZN => ATT1_n_23);
  ATT1_PM4_state2_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_15, D => ATT1_n_6, Q => FE_PHN114_ATT1_PM4_state2_0);
  ATT1_PM4_state1_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => ATT1_n_5, Q => ATT1_PM4_state1_0);
  ATT1_g817 : AOI31D0BWP7T port map(A1 => char2posx(6), A2 => char2posx(5), A3 => char2posx(7), B => char2death, ZN => ATT1_n_22);
  ATT1_g818 : INR4D0BWP7T port map(A1 => FE_PHN98_inputsp2_5, B1 => FE_OFN3_reset, B2 => ATT1_PM2_state2_0, B3 => ATT1_at2b, ZN => ATT1_n_21);
  ATT1_g819 : INR4D0BWP7T port map(A1 => inputsp2(4), B1 => ATT1_PM2_state2_1, B2 => ATT1_at2b, B3 => FE_PHN98_inputsp2_5, ZN => ATT1_n_20);
  ATT1_g820 : AOI31D0BWP7T port map(A1 => char1posx(6), A2 => char1posx(5), A3 => char1posx(7), B => char1death, ZN => ATT1_n_19);
  ATT1_g821 : AOI21D0BWP7T port map(A1 => ATT1_n_1, A2 => inputsp1(5), B => ATT1_PM2_state1_0, ZN => ATT1_n_15);
  ATT1_g822 : INR3D0BWP7T port map(A1 => inputsp1(4), B1 => ATT1_at1b, B2 => inputsp1(5), ZN => ATT1_n_14);
  ATT1_g823 : INR3D0BWP7T port map(A1 => ATT1_n_827, B1 => FE_OFN3_reset, B2 => ATT1_n_828, ZN => ATT1_n_18);
  ATT1_g824 : INR3D0BWP7T port map(A1 => ATT1_n_817, B1 => FE_OFN3_reset, B2 => ATT1_n_818, ZN => ATT1_n_17);
  ATT1_g825 : AN2D0BWP7T port map(A1 => ATT1_PM2_state2_0, A2 => ATT1_n_7, Z => ATT1_n_16);
  ATT1_g826 : INVD1BWP7T port map(I => FE_PHN146_ATT1_n_12, ZN => ATT1_n_13);
  ATT1_g827 : INVD1BWP7T port map(I => ATT1_n_10, ZN => ATT1_n_11);
  ATT1_g828 : NR4D0BWP7T port map(A1 => char2posx(2), A2 => char2posx(3), A3 => char2posx(1), A4 => char2posx(0), ZN => ATT1_n_9);
  ATT1_g829 : NR4D0BWP7T port map(A1 => char1posx(2), A2 => char1posx(3), A3 => char1posx(1), A4 => char1posx(0), ZN => ATT1_n_8);
  ATT1_g830 : IND3D1BWP7T port map(A1 => ATT1_PM2_state1_0, B1 => FE_DBTN14_reset, B2 => FE_PHN116_ATT1_PM2_state1_1, ZN => ATT1_n_12);
  ATT1_g831 : IND3D1BWP7T port map(A1 => ATT1_PM2_state2_0, B1 => FE_DBTN14_reset, B2 => ATT1_PM2_state2_1, ZN => ATT1_n_10);
  ATT1_g833 : IND2D1BWP7T port map(A1 => ATT1_PM4_state2_1, B1 => ATT1_PM4_state2_0, ZN => ATT1_n_6);
  ATT1_g834 : AN2D1BWP7T port map(A1 => Vsync, A2 => FE_DBTN14_reset, Z => ATT1_n_7);
  ATT1_g835 : IND2D1BWP7T port map(A1 => ATT1_PM4_state1_1, B1 => ATT1_PM4_state1_0, ZN => FE_PHN48_ATT1_n_5);
  ATT1_g836 : ND2D0BWP7T port map(A1 => char1posx(5), A2 => char1posx(6), ZN => ATT1_n_4);
  ATT1_g837 : ND2D0BWP7T port map(A1 => char2posx(5), A2 => char2posx(6), ZN => ATT1_n_3);
  ATT1_g14164 : INR3D0BWP7T port map(A1 => ATT1_PM2_state2_0, B1 => ATT1_PM2_state2_1, B2 => FE_OFN3_reset, ZN => ATT1_n_0);
  ATT1_PM3_state1_reg_1 : DFD1BWP7T port map(CP => CTS_17, D => ATT1_n_24, Q => ATT1_PM3_state1_1, QN => ATT1_n_62);
  ATT1_PM3_state2_reg_1 : DFD1BWP7T port map(CP => CTS_17, D => ATT1_n_23, Q => ATT1_PM3_state2_1, QN => ATT1_n_47);
  ATT1_PM3_state2_reg_0 : DFKCND1BWP7T port map(CN => ATT1_n_17, CP => CTS_17, D => ATT1_at1a, Q => ATT1_PM3_state2_0, QN => ATT1_n_44);
  ATT1_PM3_state1_reg_0 : DFKCND1BWP7T port map(CN => ATT1_n_18, CP => CTS_17, D => ATT1_at2a, Q => ATT1_PM3_state1_0, QN => ATT1_n_43);
  ATT1_PM2_state1_reg_2 : DFD1BWP7T port map(CP => CTS_16, D => FE_PHN156_ATT1_n_26, Q => ATT1_at1b, QN => ATT1_n_1);
  TL04_g3 : INVD5BWP7T port map(I => TL04_n_38, ZN => controller_clk);
  TL04_g4 : INVD0BWP7T port map(I => p2_controller, ZN => TL04_n_31);
  TL04_g5 : INVD0BWP7T port map(I => p1_controller, ZN => TL04_n_30);
  TL04_desrlzr_buttons_signal_p1_reg_7 : DFKCNQD1BWP7T port map(CN => TL04_deserializer_out_p1(6), CP => TL04_des_clk_buffered, D => TL04_n_36, Q => TL04_deserializer_out_p1(7));
  TL04_desrlzr_buttons_signal_p2_reg_7 : DFKCNQD1BWP7T port map(CN => TL04_deserializer_out_p2(6), CP => TL04_des_clk_buffered, D => TL04_n_36, Q => TL04_deserializer_out_p2(7));
  TL04_desrlzr_buttons_signal_p2_reg_6 : DFKCNQD1BWP7T port map(CN => TL04_deserializer_out_p2(5), CP => TL04_des_clk_buffered, D => TL04_n_36, Q => TL04_deserializer_out_p2(6));
  TL04_desrlzr_buttons_signal_p1_reg_6 : DFKCNQD1BWP7T port map(CN => TL04_deserializer_out_p1(5), CP => TL04_des_clk_buffered, D => TL04_n_36, Q => TL04_deserializer_out_p1(6));
  TL04_desrlzr_buttons_signal_p2_reg_5 : DFKCNQD1BWP7T port map(CN => TL04_deserializer_out_p2(4), CP => TL04_des_clk_buffered, D => TL04_n_36, Q => TL04_deserializer_out_p2(5));
  TL04_desrlzr_buttons_signal_p1_reg_5 : DFKCNQD1BWP7T port map(CN => TL04_deserializer_out_p1(4), CP => TL04_des_clk_buffered, D => TL04_n_36, Q => TL04_deserializer_out_p1(5));
  TL04_desrlzr_buttons_signal_p2_reg_4 : DFKCNQD1BWP7T port map(CN => TL04_deserializer_out_p2(3), CP => TL04_des_clk_buffered, D => TL04_n_36, Q => TL04_deserializer_out_p2(4));
  TL04_desrlzr_buttons_signal_p1_reg_4 : DFKCNQD1BWP7T port map(CN => TL04_deserializer_out_p1(3), CP => TL04_des_clk_buffered, D => TL04_n_36, Q => TL04_deserializer_out_p1(4));
  TL04_desrlzr_buttons_signal_p2_reg_3 : DFKCNQD1BWP7T port map(CN => TL04_deserializer_out_p2(2), CP => TL04_des_clk_buffered, D => TL04_n_36, Q => TL04_deserializer_out_p2(3));
  TL04_desrlzr_buttons_signal_p1_reg_3 : DFKCNQD1BWP7T port map(CN => TL04_deserializer_out_p1(2), CP => TL04_des_clk_buffered, D => TL04_n_36, Q => TL04_deserializer_out_p1(3));
  TL04_desrlzr_buttons_signal_p2_reg_2 : DFKCNQD1BWP7T port map(CN => TL04_deserializer_out_p2(1), CP => TL04_des_clk_buffered, D => TL04_n_36, Q => TL04_deserializer_out_p2(2));
  TL04_desrlzr_buttons_signal_p1_reg_2 : DFKCNQD1BWP7T port map(CN => TL04_deserializer_out_p1(1), CP => TL04_des_clk_buffered, D => TL04_n_36, Q => TL04_deserializer_out_p1(2));
  TL04_desrlzr_buttons_signal_p1_reg_1 : DFKCNQD1BWP7T port map(CN => TL04_deserializer_out_p1(0), CP => TL04_des_clk_buffered, D => TL04_n_36, Q => TL04_deserializer_out_p1(1));
  TL04_desrlzr_buttons_signal_p2_reg_1 : DFKCNQD1BWP7T port map(CN => TL04_deserializer_out_p2(0), CP => TL04_des_clk_buffered, D => TL04_n_36, Q => TL04_deserializer_out_p2(1));
  TL04_desrlzr_buttons_signal_p1_reg_0 : DFKCNQD1BWP7T port map(CN => TL04_n_30, CP => TL04_des_clk_buffered, D => TL04_n_36, Q => TL04_deserializer_out_p1(0));
  TL04_desrlzr_buttons_signal_p2_reg_0 : DFKCNQD1BWP7T port map(CN => TL04_n_31, CP => TL04_des_clk_buffered, D => TL04_n_36, Q => TL04_deserializer_out_p2(0));
  TL04_g38 : ND2D0BWP7T port map(A1 => TL04_n_36, A2 => TL04_n_33, ZN => TL04_count_reset);
  TL04_des_buffer_tmp_reg : DFQD0BWP7T port map(CP => CTS_16, D => TL04_n_28, Q => TL04_des_clk_buffered);
  TL04_g40 : OR2D1BWP7T port map(A1 => TL04_n_37, A2 => FE_PHN113_TL04_driver_state_0, Z => TL04_n_36);
  TL04_g41 : CKAN2D8BWP7T port map(A1 => TL04_n_29, A2 => FE_PHN113_TL04_driver_state_0, Z => controller_latch);
  TL04_g42 : ND4D0BWP7T port map(A1 => TL04_count(3), A2 => TL04_count(2), A3 => TL04_count(1), A4 => TL04_count(0), ZN => TL04_n_33);
  TL04_g43 : OR2D1BWP7T port map(A1 => TL04_jump_p2_state_1, A2 => TL04_jump_p2_state_0, Z => inputsp2(2));
  TL04_g44 : ND2D1BWP7T port map(A1 => TL04_driver_state_1, A2 => FE_PHN113_TL04_driver_state_0, ZN => TL04_n_38);
  TL04_g45 : INVD0BWP7T port map(I => TL04_n_29, ZN => TL04_n_37);
  TL04_g46 : NR2XD0BWP7T port map(A1 => FE_PHN113_TL04_driver_state_0, A2 => FE_OFN3_reset, ZN => TL04_n_28);
  TL04_g47 : OR2D1BWP7T port map(A1 => TL04_jump_p1_state_1, A2 => TL04_jump_p1_state_0, Z => inputsp1(2));
  TL04_g48 : NR2XD0BWP7T port map(A1 => TL04_driver_state_1, A2 => TL04_driver_state_2, ZN => TL04_n_29);
  TL04_driver_pulse_count_reg_2 : DFKCNQD1BWP7T port map(CN => TL04_n_24, CP => CTS_16, D => FE_PHN125_TL04_n_27, Q => TL04_driver_pulse_count_2);
  TL04_driver_state_reg_1 : DFQD1BWP7T port map(CP => CTS_16, D => TL04_n_26, Q => FE_PHN104_TL04_driver_state_1);
  TL04_g460 : MOAI22D0BWP7T port map(A1 => TL04_driver_pulse_count_2, A2 => TL04_n_22, B1 => TL04_driver_pulse_count_2, B2 => TL04_n_22, ZN => TL04_n_27);
  TL04_driver_pulse_count_reg_1 : DFKCNQD1BWP7T port map(CN => TL04_n_24, CP => CTS_16, D => TL04_n_23, Q => TL04_driver_pulse_count_1);
  TL04_g463 : NR3D0BWP7T port map(A1 => TL04_n_19, A2 => FE_OFN3_reset, A3 => TL04_n_25, ZN => TL04_n_26);
  TL04_driver_pulse_count_reg_0 : DFKCNQD1BWP7T port map(CN => TL04_n_16, CP => CTS_16, D => TL04_n_24, Q => FE_PHN80_TL04_driver_pulse_count_0);
  TL04_g465 : OAI21D0BWP7T port map(A1 => TL04_driver_state_1, A2 => TL04_n_21, B => TL04_n_9, ZN => TL04_n_25);
  TL04_driver_state_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL04_n_20, Q => TL04_driver_state_0);
  TL04_g467 : MOAI22D0BWP7T port map(A1 => TL04_driver_pulse_count_1, A2 => TL04_n_14, B1 => TL04_driver_pulse_count_1, B2 => TL04_n_14, ZN => FE_PHN129_TL04_n_23);
  TL04_g468 : OA31D1BWP7T port map(A1 => TL04_n_33, A2 => FE_PHN89_TL04_n_0, A3 => TL04_n_17, B => FE_PHN155_TL04_n_15, Z => TL04_n_24);
  TL04_reg_buttons_p1_reg_6 : EDFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL04_deserializer_out_p1(6), E => TL04_n_7, Q => inputsp1(6));
  TL04_reg_buttons_p1_reg_3 : EDFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL04_deserializer_out_p1(3), E => TL04_n_7, Q => inputsp1(3));
  TL04_reg_buttons_p1_reg_4 : EDFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL04_deserializer_out_p1(4), E => TL04_n_7, Q => inputsp1(4));
  TL04_reg_buttons_p1_reg_5 : EDFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL04_deserializer_out_p1(5), E => TL04_n_7, Q => inputsp1(5));
  TL04_reg_buttons_p2_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL04_deserializer_out_p2(1), E => TL04_n_7, Q => inputsp2(1));
  TL04_reg_buttons_p1_reg_7 : EDFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL04_deserializer_out_p1(7), E => TL04_n_7, Q => inputsp1(7));
  TL04_reg_buttons_p2_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL04_deserializer_out_p2(0), E => TL04_n_7, Q => inputsp2(0));
  TL04_g477 : IND2D1BWP7T port map(A1 => TL04_n_14, B1 => TL04_driver_pulse_count_1, ZN => TL04_n_22);
  TL04_reg_buttons_p2_reg_3 : EDFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL04_deserializer_out_p2(3), E => TL04_n_7, Q => inputsp2(3));
  TL04_reg_buttons_p2_reg_4 : EDFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL04_deserializer_out_p2(4), E => TL04_n_7, Q => inputsp2(4));
  TL04_reg_buttons_p2_reg_5 : EDFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL04_deserializer_out_p2(5), E => TL04_n_7, Q => inputsp2(5));
  TL04_reg_buttons_p2_reg_6 : EDFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL04_deserializer_out_p2(6), E => TL04_n_7, Q => inputsp2(6));
  TL04_reg_buttons_p2_reg_7 : EDFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL04_deserializer_out_p2(7), E => TL04_n_7, Q => inputsp2(7));
  TL04_reg_buttons_p1_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL04_deserializer_out_p1(0), E => TL04_n_7, Q => inputsp1(0));
  TL04_reg_buttons_p1_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL04_deserializer_out_p1(1), E => TL04_n_7, Q => inputsp1(1));
  TL04_jump_p1_state_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => FE_PHN64_TL04_n_12, Q => TL04_jump_p1_state_1);
  TL04_g489 : INR2XD0BWP7T port map(A1 => TL04_n_17, B1 => TL04_n_33, ZN => TL04_n_21);
  TL04_g490 : AO211D0BWP7T port map(A1 => FE_PHN113_TL04_driver_state_0, A2 => TL04_n_33, B => TL04_n_19, C => TL04_n_6, Z => TL04_n_20);
  TL04_jump_p2_state_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_15, D => FE_PHN65_TL04_n_10, Q => TL04_jump_p2_state_1);
  TL04_g492 : AN2D0BWP7T port map(A1 => FE_PHN170_TL04_n_15, A2 => TL04_n_37, Z => TL04_n_18);
  TL04_g493 : OAI21D0BWP7T port map(A1 => TL04_n_8, A2 => FE_PHN89_TL04_n_0, B => TL04_n_36, ZN => TL04_n_19);
  TL04_g494 : MOAI22D0BWP7T port map(A1 => FE_PHN173_TL04_driver_pulse_count_0, A2 => TL04_n_9, B1 => TL04_driver_pulse_count_0, B2 => TL04_n_9, ZN => TL04_n_16);
  TL04_g495 : IND4D0BWP7T port map(A1 => FE_PHN113_TL04_driver_state_0, B1 => TL04_driver_pulse_count_2, B2 => TL04_driver_pulse_count_0, B3 => TL04_driver_pulse_count_1, ZN => TL04_n_17);
  TL04_g496 : MOAI22D0BWP7T port map(A1 => inputsp1(2), A2 => TL04_n_1, B1 => TL04_jump_p1_state_0, B2 => Vsync, ZN => TL04_n_13);
  TL04_g497 : AOI21D0BWP7T port map(A1 => TL04_driver_state_2, A2 => TL04_driver_state_1, B => FE_OFN3_reset, ZN => TL04_n_15);
  TL04_g498 : IND2D1BWP7T port map(A1 => TL04_n_9, B1 => TL04_driver_pulse_count_0, ZN => TL04_n_14);
  TL04_g499 : MOAI22D0BWP7T port map(A1 => TL04_n_2, A2 => Vsync, B1 => TL04_jump_p1_state_1, B2 => TL04_jump_button_p1, ZN => TL04_n_12);
  TL04_g500 : MOAI22D0BWP7T port map(A1 => inputsp2(2), A2 => TL04_n_4, B1 => TL04_jump_p2_state_0, B2 => Vsync, ZN => TL04_n_11);
  TL04_g501 : MOAI22D0BWP7T port map(A1 => TL04_n_5, A2 => Vsync, B1 => TL04_jump_p2_state_1, B2 => TL04_jump_button_p2, ZN => TL04_n_10);
  TL04_g502 : NR2XD0BWP7T port map(A1 => FE_PHN113_TL04_driver_state_0, A2 => TL04_driver_state_1, ZN => TL04_n_8);
  TL04_g503 : OR2D1BWP7T port map(A1 => TL04_n_38, A2 => TL04_n_33, Z => TL04_n_9);
  TL04_g504 : NR2D0BWP7T port map(A1 => FE_PHN113_TL04_driver_state_0, A2 => TL04_n_33, ZN => TL04_n_6);
  TL04_g505 : AN2D1BWP7T port map(A1 => TL04_driver_state_2, A2 => FE_PHN113_TL04_driver_state_0, Z => TL04_n_7);
  TL04_jump_p2_state_reg_0 : DFKCND1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_15, D => FE_PHN78_TL04_n_11, Q => TL04_jump_p2_state_0, QN => TL04_n_5);
  TL04_reg_buttons_p2_reg_2 : EDFKCND1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL04_deserializer_out_p2(2), E => TL04_n_7, Q => TL04_jump_button_p2, QN => TL04_n_4);
  TL04_jump_p1_state_reg_0 : DFKCND1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => FE_PHN74_TL04_n_13, Q => TL04_jump_p1_state_0, QN => TL04_n_2);
  TL04_reg_buttons_p1_reg_2 : EDFKCND1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL04_deserializer_out_p1(2), E => TL04_n_7, Q => TL04_jump_button_p1, QN => TL04_n_1);
  TL04_driver_state_reg_2 : DFKCND1BWP7T port map(CN => TL04_n_25, CP => CTS_16, D => TL04_n_18, Q => TL04_driver_state_2, QN => TL04_n_0);
  TL02_PHS1_knockback_mul_35_64_g1683 : OAI31D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_97, A2 => TL02_PHS1_knockback_mul_35_64_n_122, A3 => TL02_PHS1_knockback_mul_35_64_n_171, B => TL02_PHS1_knockback_mul_35_64_n_173, ZN => TL02_n_454);
  TL02_PHS1_knockback_mul_35_64_g1684 : AO31D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_171, A2 => TL02_PHS1_knockback_mul_35_64_n_122, A3 => TL02_PHS1_knockback_mul_35_64_n_97, B => TL02_PHS1_knockback_mul_35_64_n_96, Z => TL02_PHS1_knockback_mul_35_64_n_173);
  TL02_PHS1_knockback_mul_35_64_g1685 : MOAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_171, A2 => TL02_PHS1_knockback_mul_35_64_n_129, B1 => TL02_PHS1_knockback_mul_35_64_n_171, B2 => TL02_PHS1_knockback_mul_35_64_n_129, ZN => TL02_n_456);
  TL02_PHS1_knockback_mul_35_64_g1686 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_136, B => TL02_PHS1_knockback_mul_35_64_n_121, CI => TL02_PHS1_knockback_mul_35_64_n_168, CO => TL02_PHS1_knockback_mul_35_64_n_171, S => TL02_n_457);
  TL02_PHS1_knockback_mul_35_64_g1687 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_141, B => TL02_PHS1_knockback_mul_35_64_n_137, CI => TL02_PHS1_knockback_mul_35_64_n_166, CO => TL02_PHS1_knockback_mul_35_64_n_168, S => TL02_n_458);
  TL02_PHS1_knockback_mul_35_64_g1688 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_142, B => TL02_PHS1_knockback_mul_35_64_n_148, CI => TL02_PHS1_knockback_mul_35_64_n_164, CO => TL02_PHS1_knockback_mul_35_64_n_166, S => TL02_n_459);
  TL02_PHS1_knockback_mul_35_64_g1689 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_149, B => TL02_PHS1_knockback_mul_35_64_n_156, CI => TL02_PHS1_knockback_mul_35_64_n_162, CO => TL02_PHS1_knockback_mul_35_64_n_164, S => TL02_n_460);
  TL02_PHS1_knockback_mul_35_64_g1690 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_157, B => TL02_PHS1_knockback_mul_35_64_n_153, CI => TL02_PHS1_knockback_mul_35_64_n_160, CO => TL02_PHS1_knockback_mul_35_64_n_162, S => TL02_n_461);
  TL02_PHS1_knockback_mul_35_64_g1691 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_154, B => TL02_PHS1_knockback_mul_35_64_n_151, CI => TL02_PHS1_knockback_mul_35_64_n_158, CO => TL02_PHS1_knockback_mul_35_64_n_160, S => TL02_n_462);
  TL02_PHS1_knockback_mul_35_64_g1692 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_152, B => TL02_PHS1_knockback_mul_35_64_n_144, CI => TL02_PHS1_knockback_mul_35_64_n_155, CO => TL02_PHS1_knockback_mul_35_64_n_158, S => TL02_n_463);
  TL02_PHS1_knockback_mul_35_64_g1693 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_146, B => TL02_PHS1_knockback_mul_35_64_n_105, CI => TL02_PHS1_knockback_mul_35_64_n_124, CO => TL02_PHS1_knockback_mul_35_64_n_156, S => TL02_PHS1_knockback_mul_35_64_n_157);
  TL02_PHS1_knockback_mul_35_64_g1694 : MAOI222D1BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_150, B => TL02_PHS1_knockback_mul_35_64_n_143, C => TL02_PHS1_knockback_mul_35_64_n_134, ZN => TL02_PHS1_knockback_mul_35_64_n_155);
  TL02_PHS1_knockback_mul_35_64_g1695 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_138, B => TL02_PHS1_knockback_mul_35_64_n_109, CI => TL02_PHS1_knockback_mul_35_64_n_147, CO => TL02_PHS1_knockback_mul_35_64_n_153, S => TL02_PHS1_knockback_mul_35_64_n_154);
  TL02_PHS1_knockback_mul_35_64_g1696 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_116, B => TL02_PHS1_knockback_mul_35_64_n_70, CI => TL02_PHS1_knockback_mul_35_64_n_139, CO => TL02_PHS1_knockback_mul_35_64_n_151, S => TL02_PHS1_knockback_mul_35_64_n_152);
  TL02_PHS1_knockback_mul_35_64_g1697 : MAOI222D1BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_145, B => TL02_PHS1_knockback_mul_35_64_n_199, C => TL02_PHS1_knockback_mul_35_64_n_117, ZN => TL02_PHS1_knockback_mul_35_64_n_150);
  TL02_PHS1_knockback_mul_35_64_g1698 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_123, B => TL02_PHS1_knockback_mul_35_64_n_100, CI => TL02_PHS1_knockback_mul_35_64_n_126, CO => TL02_PHS1_knockback_mul_35_64_n_148, S => TL02_PHS1_knockback_mul_35_64_n_149);
  TL02_PHS1_knockback_mul_35_64_g1699 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_67, B => TL02_PHS1_knockback_mul_35_64_n_127, CI => TL02_PHS1_knockback_mul_35_64_n_66, CO => TL02_PHS1_knockback_mul_35_64_n_146, S => TL02_PHS1_knockback_mul_35_64_n_147);
  TL02_PHS1_knockback_mul_35_64_g1700 : MAOI222D1BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_130, B => TL02_PHS1_knockback_mul_35_64_n_135, C => TL02_PHS1_knockback_mul_35_64_n_110, ZN => TL02_PHS1_knockback_mul_35_64_n_145);
  TL02_PHS1_knockback_mul_35_64_g1701 : MAOI222D1BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_131, B => TL02_PHS1_knockback_mul_35_64_n_63, C => TL02_PHS1_knockback_mul_35_64_n_111, ZN => TL02_PHS1_knockback_mul_35_64_n_144);
  TL02_PHS1_knockback_mul_35_64_g1702 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_132, A2 => TL02_PHS1_knockback_mul_35_64_n_131, B1 => TL02_PHS1_knockback_mul_35_64_n_132, B2 => TL02_PHS1_knockback_mul_35_64_n_131, ZN => TL02_PHS1_knockback_mul_35_64_n_143);
  TL02_PHS1_knockback_mul_35_64_g1703 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_125, B => TL02_PHS1_knockback_mul_35_64_n_71, CI => TL02_PHS1_knockback_mul_35_64_n_120, CO => TL02_PHS1_knockback_mul_35_64_n_141, S => TL02_PHS1_knockback_mul_35_64_n_142);
  TL02_PHS1_knockback_mul_35_64_g1705 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_128, B => TL02_PHS1_knockback_mul_35_64_n_83, CI => TL02_PHS1_knockback_mul_35_64_n_64, CO => TL02_PHS1_knockback_mul_35_64_n_138, S => TL02_PHS1_knockback_mul_35_64_n_139);
  TL02_PHS1_knockback_mul_35_64_g1706 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_68, B => TL02_PHS1_knockback_mul_35_64_n_91, CI => TL02_PHS1_knockback_mul_35_64_n_119, CO => TL02_PHS1_knockback_mul_35_64_n_136, S => TL02_PHS1_knockback_mul_35_64_n_137);
  TL02_PHS1_knockback_mul_35_64_g1707 : MAOI222D1BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_112, B => TL02_PHS1_knockback_mul_35_64_n_201, C => TL02_PHS1_knockback_mul_35_64_n_58, ZN => TL02_PHS1_knockback_mul_35_64_n_135);
  TL02_PHS1_knockback_mul_35_64_g1708 : MAOI222D1BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_60, B => TL02_PHS1_knockback_mul_35_64_n_114, C => TL02_PHS1_knockback_mul_35_64_n_77, ZN => TL02_PHS1_knockback_mul_35_64_n_134);
  TL02_PHS1_knockback_mul_35_64_g1710 : CKXOR2D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_63, A2 => TL02_PHS1_knockback_mul_35_64_n_111, Z => TL02_PHS1_knockback_mul_35_64_n_132);
  TL02_PHS1_knockback_mul_35_64_g1711 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_74, A2 => TL02_PHS1_knockback_mul_35_64_n_115, B1 => TL02_PHS1_knockback_mul_35_64_n_74, B2 => TL02_PHS1_knockback_mul_35_64_n_115, ZN => TL02_PHS1_knockback_mul_35_64_n_131);
  TL02_PHS1_knockback_mul_35_64_g1712 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_59, A2 => TL02_PHS1_knockback_mul_35_64_n_113, B1 => TL02_PHS1_knockback_mul_35_64_n_59, B2 => TL02_PHS1_knockback_mul_35_64_n_113, ZN => TL02_PHS1_knockback_mul_35_64_n_130);
  TL02_PHS1_knockback_mul_35_64_g1713 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_122, A2 => TL02_PHS1_knockback_mul_35_64_n_97, B1 => TL02_PHS1_knockback_mul_35_64_n_122, B2 => TL02_PHS1_knockback_mul_35_64_n_97, ZN => TL02_PHS1_knockback_mul_35_64_n_129);
  TL02_PHS1_knockback_mul_35_64_g1714 : HA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_102, B => TL02_PHS1_knockback_mul_35_64_n_73, CO => TL02_PHS1_knockback_mul_35_64_n_127, S => TL02_PHS1_knockback_mul_35_64_n_128);
  TL02_PHS1_knockback_mul_35_64_g1715 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_82, B => TL02_PHS1_knockback_mul_35_64_n_89, CI => TL02_PHS1_knockback_mul_35_64_n_86, CO => TL02_PHS1_knockback_mul_35_64_n_125, S => TL02_PHS1_knockback_mul_35_64_n_126);
  TL02_PHS1_knockback_mul_35_64_g1716 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_84, B => TL02_PHS1_knockback_mul_35_64_n_108, CI => TL02_PHS1_knockback_mul_35_64_n_65, CO => TL02_PHS1_knockback_mul_35_64_n_123, S => TL02_PHS1_knockback_mul_35_64_n_124);
  TL02_PHS1_knockback_mul_35_64_g1717 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_92, B => TL02_PHS1_knockback_mul_35_64_n_93, CI => TL02_PHS1_knockback_mul_35_64_n_69, CO => TL02_PHS1_knockback_mul_35_64_n_122, S => TL02_PHS1_knockback_mul_35_64_n_121);
  TL02_PHS1_knockback_mul_35_64_g1718 : FA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_90, B => TL02_PHS1_knockback_mul_35_64_n_94, CI => TL02_PHS1_knockback_mul_35_64_n_85, CO => TL02_PHS1_knockback_mul_35_64_n_119, S => TL02_PHS1_knockback_mul_35_64_n_120);
  TL02_PHS1_knockback_mul_35_64_g1720 : MAOI222D1BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_59, B => TL02_PHS1_knockback_mul_35_64_n_76, C => TL02_PHS1_knockback_mul_35_64_n_104, ZN => TL02_PHS1_knockback_mul_35_64_n_117);
  TL02_PHS1_knockback_mul_35_64_g1721 : MAOI222D1BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_75, B => TL02_PHS1_knockback_mul_35_64_n_78, C => TL02_PHS1_knockback_mul_35_64_n_103, ZN => TL02_PHS1_knockback_mul_35_64_n_116);
  TL02_PHS1_knockback_mul_35_64_g1722 : XNR2D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_78, A2 => TL02_PHS1_knockback_mul_35_64_n_103, ZN => TL02_PHS1_knockback_mul_35_64_n_115);
  TL02_PHS1_knockback_mul_35_64_g1723 : MOAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_79, A2 => TL02_PHS1_knockback_mul_35_64_n_101, B1 => TL02_PHS1_knockback_mul_35_64_n_79, B2 => TL02_PHS1_knockback_mul_35_64_n_101, ZN => TL02_PHS1_knockback_mul_35_64_n_114);
  TL02_PHS1_knockback_mul_35_64_g1724 : CKXOR2D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_76, A2 => TL02_PHS1_knockback_mul_35_64_n_104, Z => TL02_PHS1_knockback_mul_35_64_n_113);
  TL02_PHS1_knockback_mul_35_64_g1725 : MOAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_80, A2 => TL02_PHS1_knockback_mul_35_64_n_107, B1 => TL02_PHS1_knockback_mul_35_64_n_80, B2 => TL02_PHS1_knockback_mul_35_64_n_107, ZN => TL02_PHS1_knockback_mul_35_64_n_112);
  TL02_PHS1_knockback_mul_35_64_g1726 : IND2D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_79, B1 => TL02_PHS1_knockback_mul_35_64_n_101, ZN => TL02_PHS1_knockback_mul_35_64_n_111);
  TL02_PHS1_knockback_mul_35_64_g1727 : IND2D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_80, B1 => TL02_PHS1_knockback_mul_35_64_n_107, ZN => TL02_PHS1_knockback_mul_35_64_n_110);
  TL02_PHS1_knockback_mul_35_64_g1728 : HA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_62, B => TL02_PHS1_knockback_mul_35_64_n_72, CO => TL02_PHS1_knockback_mul_35_64_n_108, S => TL02_PHS1_knockback_mul_35_64_n_109);
  TL02_PHS1_knockback_mul_35_64_g1729 : HA1D0BWP7T port map(A => TL02_PHS1_knockback_mul_35_64_n_95, B => TL02_PHS1_knockback_mul_35_64_n_87, CO => TL02_PHS1_knockback_mul_35_64_n_107, S => TL02_PHS1_knockback_mul_35_64_n_106);
  TL02_PHS1_knockback_mul_35_64_g1730 : OAI21D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_81, A2 => TL02_n_444, B => TL02_PHS1_knockback_mul_35_64_n_100, ZN => TL02_PHS1_knockback_mul_35_64_n_105);
  TL02_PHS1_knockback_mul_35_64_g1731 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_99, A2 => TL02_PHS1_knockback_mul_35_64_n_93, B1 => TL02_PHS1_knockback_mul_35_64_n_99, B2 => TL02_PHS1_knockback_mul_35_64_n_93, ZN => TL02_PHS1_knockback_mul_35_64_n_104);
  TL02_PHS1_knockback_mul_35_64_g1732 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_98, A2 => TL02_PHS1_knockback_mul_35_64_n_96, B1 => TL02_PHS1_knockback_mul_35_64_n_98, B2 => TL02_PHS1_knockback_mul_35_64_n_96, ZN => TL02_PHS1_knockback_mul_35_64_n_103);
  TL02_PHS1_knockback_mul_35_64_g1733 : INR2XD0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_98, B1 => TL02_PHS1_knockback_mul_35_64_n_96, ZN => TL02_PHS1_knockback_mul_35_64_n_102);
  TL02_PHS1_knockback_mul_35_64_g1734 : INR2D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_99, B1 => TL02_PHS1_knockback_mul_35_64_n_93, ZN => TL02_PHS1_knockback_mul_35_64_n_101);
  TL02_PHS1_knockback_mul_35_64_g1735 : ND2D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_81, A2 => TL02_n_444, ZN => TL02_PHS1_knockback_mul_35_64_n_100);
  TL02_PHS1_knockback_mul_35_64_g1736 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_35_64_n_94, ZN => TL02_PHS1_knockback_mul_35_64_n_95);
  TL02_PHS1_knockback_mul_35_64_g1737 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_35_64_n_91, ZN => TL02_PHS1_knockback_mul_35_64_n_92);
  TL02_PHS1_knockback_mul_35_64_g1738 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_35_64_n_89, ZN => TL02_PHS1_knockback_mul_35_64_n_90);
  TL02_PHS1_knockback_mul_35_64_g1740 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_55, A2 => TL02_PHS1_knockback_mul_35_64_n_3, B1 => TL02_PHS1_knockback_mul_35_64_n_49, B2 => TL02_PHS1_knockback_mul_35_64_n_34, ZN => TL02_PHS1_knockback_mul_35_64_n_99);
  TL02_PHS1_knockback_mul_35_64_g1741 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_51, A2 => TL02_PHS1_knockback_mul_35_64_n_4, B1 => TL02_PHS1_knockback_mul_35_64_n_45, B2 => TL02_PHS1_knockback_mul_35_64_n_33, ZN => TL02_PHS1_knockback_mul_35_64_n_98);
  TL02_PHS1_knockback_mul_35_64_g1742 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_53, A2 => TL02_PHS1_knockback_mul_35_64_n_1, B1 => TL02_PHS1_knockback_mul_35_64_n_48, B2 => TL02_PHS1_knockback_mul_35_64_n_36, ZN => TL02_PHS1_knockback_mul_35_64_n_87);
  TL02_PHS1_knockback_mul_35_64_g1743 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_23, A2 => TL02_PHS1_knockback_mul_35_64_n_55, B1 => TL02_PHS1_knockback_mul_35_64_n_40, B2 => TL02_PHS1_knockback_mul_35_64_n_34, ZN => TL02_PHS1_knockback_mul_35_64_n_86);
  TL02_PHS1_knockback_mul_35_64_g1744 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_40, A2 => TL02_PHS1_knockback_mul_35_64_n_55, B1 => TL02_PHS1_knockback_mul_35_64_n_43, B2 => TL02_PHS1_knockback_mul_35_64_n_34, ZN => TL02_PHS1_knockback_mul_35_64_n_85);
  TL02_PHS1_knockback_mul_35_64_g1745 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_47, A2 => TL02_PHS1_knockback_mul_35_64_n_53, B1 => TL02_PHS1_knockback_mul_35_64_n_24, B2 => TL02_PHS1_knockback_mul_35_64_n_36, ZN => TL02_PHS1_knockback_mul_35_64_n_84);
  TL02_PHS1_knockback_mul_35_64_g1746 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_20, A2 => TL02_PHS1_knockback_mul_35_64_n_51, B1 => TL02_PHS1_knockback_mul_35_64_n_33, B2 => TL02_PHS1_knockback_mul_35_64_n_4, ZN => TL02_PHS1_knockback_mul_35_64_n_97);
  TL02_PHS1_knockback_mul_35_64_g1747 : OAI21D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_52, A2 => TL02_PHS1_knockback_mul_35_64_n_32, B => TL02_n_438, ZN => TL02_PHS1_knockback_mul_35_64_n_96);
  TL02_PHS1_knockback_mul_35_64_g1748 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_38, A2 => TL02_PHS1_knockback_mul_35_64_n_55, B1 => TL02_PHS1_knockback_mul_35_64_n_42, B2 => TL02_PHS1_knockback_mul_35_64_n_34, ZN => TL02_PHS1_knockback_mul_35_64_n_83);
  TL02_PHS1_knockback_mul_35_64_g1749 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_28, A2 => TL02_PHS1_knockback_mul_35_64_n_51, B1 => TL02_PHS1_knockback_mul_35_64_n_15, B2 => TL02_PHS1_knockback_mul_35_64_n_33, ZN => TL02_PHS1_knockback_mul_35_64_n_82);
  TL02_PHS1_knockback_mul_35_64_g1750 : OAI21D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_54, A2 => TL02_PHS1_knockback_mul_35_64_n_37, B => TL02_n_442, ZN => TL02_PHS1_knockback_mul_35_64_n_94);
  TL02_PHS1_knockback_mul_35_64_g1751 : OAI21D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_56, A2 => TL02_PHS1_knockback_mul_35_64_n_35, B => TL02_n_440, ZN => TL02_PHS1_knockback_mul_35_64_n_93);
  TL02_PHS1_knockback_mul_35_64_g1752 : AOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_44, A2 => TL02_PHS1_knockback_mul_35_64_n_56, B1 => TL02_PHS1_knockback_mul_35_64_n_35, B2 => TL02_n_440, ZN => TL02_PHS1_knockback_mul_35_64_n_91);
  TL02_PHS1_knockback_mul_35_64_g1753 : AOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_25, A2 => TL02_PHS1_knockback_mul_35_64_n_54, B1 => TL02_PHS1_knockback_mul_35_64_n_37, B2 => TL02_n_442, ZN => TL02_PHS1_knockback_mul_35_64_n_89);
  TL02_PHS1_knockback_mul_35_64_g1754 : INVD1BWP7T port map(I => TL02_PHS1_knockback_mul_35_64_n_74, ZN => TL02_PHS1_knockback_mul_35_64_n_75);
  TL02_PHS1_knockback_mul_35_64_g1755 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_18, A2 => TL02_PHS1_knockback_mul_35_64_n_52, B1 => TL02_PHS1_knockback_mul_35_64_n_28, B2 => TL02_PHS1_knockback_mul_35_64_n_33, ZN => TL02_PHS1_knockback_mul_35_64_n_81);
  TL02_PHS1_knockback_mul_35_64_g1756 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_45, A2 => TL02_PHS1_knockback_mul_35_64_n_51, B1 => TL02_PHS1_knockback_mul_35_64_n_14, B2 => TL02_PHS1_knockback_mul_35_64_n_33, ZN => TL02_PHS1_knockback_mul_35_64_n_73);
  TL02_PHS1_knockback_mul_35_64_g1757 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_16, A2 => TL02_PHS1_knockback_mul_35_64_n_37, B1 => TL02_PHS1_knockback_mul_35_64_n_48, B2 => TL02_PHS1_knockback_mul_35_64_n_53, ZN => TL02_PHS1_knockback_mul_35_64_n_80);
  TL02_PHS1_knockback_mul_35_64_g1758 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_22, A2 => TL02_PHS1_knockback_mul_35_64_n_35, B1 => TL02_PHS1_knockback_mul_35_64_n_49, B2 => TL02_PHS1_knockback_mul_35_64_n_55, ZN => TL02_PHS1_knockback_mul_35_64_n_79);
  TL02_PHS1_knockback_mul_35_64_g1759 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_14, A2 => TL02_PHS1_knockback_mul_35_64_n_51, B1 => TL02_PHS1_knockback_mul_35_64_n_17, B2 => TL02_PHS1_knockback_mul_35_64_n_33, ZN => TL02_PHS1_knockback_mul_35_64_n_72);
  TL02_PHS1_knockback_mul_35_64_g1760 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_15, A2 => TL02_PHS1_knockback_mul_35_64_n_51, B1 => TL02_PHS1_knockback_mul_35_64_n_21, B2 => TL02_PHS1_knockback_mul_35_64_n_33, ZN => TL02_PHS1_knockback_mul_35_64_n_71);
  TL02_PHS1_knockback_mul_35_64_g1761 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_41, A2 => TL02_PHS1_knockback_mul_35_64_n_53, B1 => TL02_PHS1_knockback_mul_35_64_n_46, B2 => TL02_PHS1_knockback_mul_35_64_n_36, ZN => TL02_PHS1_knockback_mul_35_64_n_70);
  TL02_PHS1_knockback_mul_35_64_g1762 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_19, A2 => TL02_PHS1_knockback_mul_35_64_n_51, B1 => TL02_PHS1_knockback_mul_35_64_n_20, B2 => TL02_PHS1_knockback_mul_35_64_n_33, ZN => TL02_PHS1_knockback_mul_35_64_n_69);
  TL02_PHS1_knockback_mul_35_64_g1763 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_22, A2 => TL02_PHS1_knockback_mul_35_64_n_56, B1 => TL02_PHS1_knockback_mul_35_64_n_38, B2 => TL02_PHS1_knockback_mul_35_64_n_34, ZN => TL02_PHS1_knockback_mul_35_64_n_78);
  TL02_PHS1_knockback_mul_35_64_g1764 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_27, A2 => TL02_PHS1_knockback_mul_35_64_n_53, B1 => TL02_PHS1_knockback_mul_35_64_n_39, B2 => TL02_PHS1_knockback_mul_35_64_n_36, ZN => TL02_PHS1_knockback_mul_35_64_n_77);
  TL02_PHS1_knockback_mul_35_64_g1765 : AOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_16, A2 => TL02_PHS1_knockback_mul_35_64_n_54, B1 => TL02_PHS1_knockback_mul_35_64_n_26, B2 => TL02_PHS1_knockback_mul_35_64_n_37, ZN => TL02_PHS1_knockback_mul_35_64_n_76);
  TL02_PHS1_knockback_mul_35_64_g1766 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_21, A2 => TL02_PHS1_knockback_mul_35_64_n_51, B1 => TL02_PHS1_knockback_mul_35_64_n_19, B2 => TL02_PHS1_knockback_mul_35_64_n_33, ZN => TL02_PHS1_knockback_mul_35_64_n_68);
  TL02_PHS1_knockback_mul_35_64_g1767 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_42, A2 => TL02_PHS1_knockback_mul_35_64_n_55, B1 => TL02_PHS1_knockback_mul_35_64_n_50, B2 => TL02_PHS1_knockback_mul_35_64_n_34, ZN => TL02_PHS1_knockback_mul_35_64_n_67);
  TL02_PHS1_knockback_mul_35_64_g1768 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_46, A2 => TL02_PHS1_knockback_mul_35_64_n_53, B1 => TL02_PHS1_knockback_mul_35_64_n_47, B2 => TL02_PHS1_knockback_mul_35_64_n_36, ZN => TL02_PHS1_knockback_mul_35_64_n_66);
  TL02_PHS1_knockback_mul_35_64_g1769 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_39, A2 => TL02_PHS1_knockback_mul_35_64_n_53, B1 => TL02_PHS1_knockback_mul_35_64_n_41, B2 => TL02_PHS1_knockback_mul_35_64_n_36, ZN => TL02_PHS1_knockback_mul_35_64_n_74);
  TL02_PHS1_knockback_mul_35_64_g1770 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_50, A2 => TL02_PHS1_knockback_mul_35_64_n_55, B1 => TL02_PHS1_knockback_mul_35_64_n_23, B2 => TL02_PHS1_knockback_mul_35_64_n_34, ZN => TL02_PHS1_knockback_mul_35_64_n_65);
  TL02_PHS1_knockback_mul_35_64_g1771 : MOAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_11, A2 => TL02_PHS1_knockback_mul_35_64_n_7, B1 => TL02_PHS1_knockback_mul_35_64_n_8, B2 => TL02_n_445, ZN => TL02_PHS1_knockback_mul_35_64_n_64);
  TL02_PHS1_knockback_mul_35_64_g1772 : OA22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_12, A2 => TL02_PHS1_knockback_mul_35_64_n_7, B1 => TL02_PHS1_knockback_mul_35_64_n_5, B2 => TL02_PHS1_knockback_mul_35_64_n_11, Z => TL02_PHS1_knockback_mul_35_64_n_63);
  TL02_PHS1_knockback_mul_35_64_g1773 : MOAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_2, A2 => TL02_PHS1_knockback_mul_35_64_n_5, B1 => TL02_PHS1_knockback_mul_35_64_n_8, B2 => TL02_PHS1_knockback_mul_35_64_n_6, ZN => TL02_PHS1_knockback_mul_35_64_n_62);
  TL02_PHS1_knockback_mul_35_64_g1775 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_10, A2 => TL02_PHS1_knockback_mul_35_64_n_7, B1 => TL02_PHS1_knockback_mul_35_64_n_12, B2 => TL02_PHS1_knockback_mul_35_64_n_5, ZN => TL02_PHS1_knockback_mul_35_64_n_60);
  TL02_PHS1_knockback_mul_35_64_g1776 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_13, A2 => TL02_PHS1_knockback_mul_35_64_n_6, B1 => TL02_PHS1_knockback_mul_35_64_n_10, B2 => TL02_PHS1_knockback_mul_35_64_n_5, ZN => TL02_PHS1_knockback_mul_35_64_n_59);
  TL02_PHS1_knockback_mul_35_64_g1777 : MOAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_9, A2 => TL02_PHS1_knockback_mul_35_64_n_7, B1 => TL02_PHS1_knockback_mul_35_64_n_13, B2 => TL02_n_445, ZN => TL02_PHS1_knockback_mul_35_64_n_58);
  TL02_PHS1_knockback_mul_35_64_g1778 : OAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_9, A2 => TL02_PHS1_knockback_mul_35_64_n_5, B1 => TL02_n_452, B2 => TL02_PHS1_knockback_mul_35_64_n_7, ZN => TL02_PHS1_knockback_mul_35_64_n_57);
  TL02_PHS1_knockback_mul_35_64_g1779 : INVD1BWP7T port map(I => TL02_PHS1_knockback_mul_35_64_n_56, ZN => TL02_PHS1_knockback_mul_35_64_n_55);
  TL02_PHS1_knockback_mul_35_64_g1780 : NR2XD0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_31, A2 => TL02_PHS1_knockback_mul_35_64_n_35, ZN => TL02_PHS1_knockback_mul_35_64_n_56);
  TL02_PHS1_knockback_mul_35_64_g1781 : INVD1BWP7T port map(I => TL02_PHS1_knockback_mul_35_64_n_54, ZN => TL02_PHS1_knockback_mul_35_64_n_53);
  TL02_PHS1_knockback_mul_35_64_g1782 : NR2XD0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_37, A2 => TL02_PHS1_knockback_mul_35_64_n_29, ZN => TL02_PHS1_knockback_mul_35_64_n_54);
  TL02_PHS1_knockback_mul_35_64_g1783 : INVD1BWP7T port map(I => TL02_PHS1_knockback_mul_35_64_n_52, ZN => TL02_PHS1_knockback_mul_35_64_n_51);
  TL02_PHS1_knockback_mul_35_64_g1784 : NR2XD0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_32, A2 => TL02_PHS1_knockback_mul_35_64_n_30, ZN => TL02_PHS1_knockback_mul_35_64_n_52);
  TL02_PHS1_knockback_mul_35_64_g1785 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_35_64_n_43, ZN => TL02_PHS1_knockback_mul_35_64_n_44);
  TL02_PHS1_knockback_mul_35_64_g1786 : INVD1BWP7T port map(I => TL02_PHS1_knockback_mul_35_64_n_37, ZN => TL02_PHS1_knockback_mul_35_64_n_36);
  TL02_PHS1_knockback_mul_35_64_g1787 : INVD1BWP7T port map(I => TL02_PHS1_knockback_mul_35_64_n_35, ZN => TL02_PHS1_knockback_mul_35_64_n_34);
  TL02_PHS1_knockback_mul_35_64_g1788 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_35_64_n_33, ZN => TL02_PHS1_knockback_mul_35_64_n_32);
  TL02_PHS1_knockback_mul_35_64_g1789 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_3, A2 => TL02_n_441, B1 => TL02_PHS1_knockback_mul_35_64_n_3, B2 => TL02_n_441, ZN => TL02_PHS1_knockback_mul_35_64_n_31);
  TL02_PHS1_knockback_mul_35_64_g1790 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_4, A2 => TL02_n_439, B1 => TL02_PHS1_knockback_mul_35_64_n_4, B2 => TL02_n_439, ZN => TL02_PHS1_knockback_mul_35_64_n_30);
  TL02_PHS1_knockback_mul_35_64_g1791 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_1, A2 => TL02_n_443, B1 => TL02_PHS1_knockback_mul_35_64_n_1, B2 => TL02_n_443, ZN => TL02_PHS1_knockback_mul_35_64_n_29);
  TL02_PHS1_knockback_mul_35_64_g1792 : MAOI22D0BWP7T port map(A1 => TL02_n_449, A2 => TL02_PHS1_knockback_mul_35_64_n_3, B1 => TL02_n_449, B2 => TL02_PHS1_knockback_mul_35_64_n_3, ZN => TL02_PHS1_knockback_mul_35_64_n_50);
  TL02_PHS1_knockback_mul_35_64_g1793 : MAOI22D0BWP7T port map(A1 => TL02_n_453, A2 => TL02_PHS1_knockback_mul_35_64_n_3, B1 => TL02_n_453, B2 => TL02_PHS1_knockback_mul_35_64_n_3, ZN => TL02_PHS1_knockback_mul_35_64_n_49);
  TL02_PHS1_knockback_mul_35_64_g1794 : MAOI22D0BWP7T port map(A1 => TL02_n_453, A2 => TL02_PHS1_knockback_mul_35_64_n_1, B1 => TL02_n_453, B2 => TL02_PHS1_knockback_mul_35_64_n_1, ZN => TL02_PHS1_knockback_mul_35_64_n_48);
  TL02_PHS1_knockback_mul_35_64_g1795 : MAOI22D0BWP7T port map(A1 => TL02_n_447, A2 => TL02_PHS1_knockback_mul_35_64_n_1, B1 => TL02_n_447, B2 => TL02_PHS1_knockback_mul_35_64_n_1, ZN => TL02_PHS1_knockback_mul_35_64_n_47);
  TL02_PHS1_knockback_mul_35_64_g1796 : MAOI22D0BWP7T port map(A1 => TL02_n_448, A2 => TL02_PHS1_knockback_mul_35_64_n_1, B1 => TL02_n_448, B2 => TL02_PHS1_knockback_mul_35_64_n_1, ZN => TL02_PHS1_knockback_mul_35_64_n_46);
  TL02_PHS1_knockback_mul_35_64_g1797 : MAOI22D0BWP7T port map(A1 => TL02_n_453, A2 => TL02_PHS1_knockback_mul_35_64_n_4, B1 => TL02_n_453, B2 => TL02_PHS1_knockback_mul_35_64_n_4, ZN => TL02_PHS1_knockback_mul_35_64_n_45);
  TL02_PHS1_knockback_mul_35_64_g1798 : MAOI22D0BWP7T port map(A1 => TL02_n_446, A2 => TL02_PHS1_knockback_mul_35_64_n_3, B1 => TL02_n_446, B2 => TL02_PHS1_knockback_mul_35_64_n_3, ZN => TL02_PHS1_knockback_mul_35_64_n_43);
  TL02_PHS1_knockback_mul_35_64_g1799 : MAOI22D0BWP7T port map(A1 => TL02_n_450, A2 => TL02_PHS1_knockback_mul_35_64_n_3, B1 => TL02_n_450, B2 => TL02_PHS1_knockback_mul_35_64_n_3, ZN => TL02_PHS1_knockback_mul_35_64_n_42);
  TL02_PHS1_knockback_mul_35_64_g1800 : MAOI22D0BWP7T port map(A1 => TL02_n_449, A2 => TL02_PHS1_knockback_mul_35_64_n_1, B1 => TL02_n_449, B2 => TL02_PHS1_knockback_mul_35_64_n_1, ZN => TL02_PHS1_knockback_mul_35_64_n_41);
  TL02_PHS1_knockback_mul_35_64_g1801 : MAOI22D0BWP7T port map(A1 => TL02_n_447, A2 => TL02_PHS1_knockback_mul_35_64_n_3, B1 => TL02_n_447, B2 => TL02_PHS1_knockback_mul_35_64_n_3, ZN => TL02_PHS1_knockback_mul_35_64_n_40);
  TL02_PHS1_knockback_mul_35_64_g1802 : MAOI22D0BWP7T port map(A1 => TL02_n_450, A2 => TL02_PHS1_knockback_mul_35_64_n_1, B1 => TL02_n_450, B2 => TL02_PHS1_knockback_mul_35_64_n_1, ZN => TL02_PHS1_knockback_mul_35_64_n_39);
  TL02_PHS1_knockback_mul_35_64_g1803 : MAOI22D0BWP7T port map(A1 => TL02_n_451, A2 => TL02_PHS1_knockback_mul_35_64_n_3, B1 => TL02_n_451, B2 => TL02_PHS1_knockback_mul_35_64_n_3, ZN => TL02_PHS1_knockback_mul_35_64_n_38);
  TL02_PHS1_knockback_mul_35_64_g1804 : MOAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_2, A2 => TL02_n_443, B1 => TL02_PHS1_knockback_mul_35_64_n_2, B2 => TL02_n_443, ZN => TL02_PHS1_knockback_mul_35_64_n_37);
  TL02_PHS1_knockback_mul_35_64_g1805 : MOAI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_1, A2 => TL02_n_441, B1 => TL02_PHS1_knockback_mul_35_64_n_1, B2 => TL02_n_441, ZN => TL02_PHS1_knockback_mul_35_64_n_35);
  TL02_PHS1_knockback_mul_35_64_g1806 : MAOI22D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_3, A2 => TL02_n_439, B1 => TL02_PHS1_knockback_mul_35_64_n_3, B2 => TL02_n_439, ZN => TL02_PHS1_knockback_mul_35_64_n_33);
  TL02_PHS1_knockback_mul_35_64_g1807 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_35_64_n_26, ZN => TL02_PHS1_knockback_mul_35_64_n_27);
  TL02_PHS1_knockback_mul_35_64_g1808 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_35_64_n_24, ZN => TL02_PHS1_knockback_mul_35_64_n_25);
  TL02_PHS1_knockback_mul_35_64_g1809 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_35_64_n_17, ZN => TL02_PHS1_knockback_mul_35_64_n_18);
  TL02_PHS1_knockback_mul_35_64_g1810 : MAOI22D0BWP7T port map(A1 => TL02_n_450, A2 => TL02_PHS1_knockback_mul_35_64_n_4, B1 => TL02_n_450, B2 => TL02_PHS1_knockback_mul_35_64_n_4, ZN => TL02_PHS1_knockback_mul_35_64_n_28);
  TL02_PHS1_knockback_mul_35_64_g1811 : MOAI22D0BWP7T port map(A1 => TL02_n_451, A2 => TL02_PHS1_knockback_mul_35_64_n_1, B1 => TL02_n_451, B2 => TL02_PHS1_knockback_mul_35_64_n_1, ZN => TL02_PHS1_knockback_mul_35_64_n_26);
  TL02_PHS1_knockback_mul_35_64_g1812 : MAOI22D0BWP7T port map(A1 => TL02_n_446, A2 => TL02_PHS1_knockback_mul_35_64_n_1, B1 => TL02_n_446, B2 => TL02_PHS1_knockback_mul_35_64_n_1, ZN => TL02_PHS1_knockback_mul_35_64_n_24);
  TL02_PHS1_knockback_mul_35_64_g1813 : MAOI22D0BWP7T port map(A1 => TL02_n_448, A2 => TL02_PHS1_knockback_mul_35_64_n_3, B1 => TL02_n_448, B2 => TL02_PHS1_knockback_mul_35_64_n_3, ZN => TL02_PHS1_knockback_mul_35_64_n_23);
  TL02_PHS1_knockback_mul_35_64_g1814 : MOAI22D0BWP7T port map(A1 => TL02_n_452, A2 => TL02_PHS1_knockback_mul_35_64_n_3, B1 => TL02_n_452, B2 => TL02_PHS1_knockback_mul_35_64_n_3, ZN => TL02_PHS1_knockback_mul_35_64_n_22);
  TL02_PHS1_knockback_mul_35_64_g1815 : MAOI22D0BWP7T port map(A1 => TL02_n_448, A2 => TL02_PHS1_knockback_mul_35_64_n_4, B1 => TL02_n_448, B2 => TL02_PHS1_knockback_mul_35_64_n_4, ZN => TL02_PHS1_knockback_mul_35_64_n_21);
  TL02_PHS1_knockback_mul_35_64_g1816 : MAOI22D0BWP7T port map(A1 => TL02_n_446, A2 => TL02_PHS1_knockback_mul_35_64_n_4, B1 => TL02_n_446, B2 => TL02_PHS1_knockback_mul_35_64_n_4, ZN => TL02_PHS1_knockback_mul_35_64_n_20);
  TL02_PHS1_knockback_mul_35_64_g1817 : MAOI22D0BWP7T port map(A1 => TL02_n_447, A2 => TL02_PHS1_knockback_mul_35_64_n_4, B1 => TL02_n_447, B2 => TL02_PHS1_knockback_mul_35_64_n_4, ZN => TL02_PHS1_knockback_mul_35_64_n_19);
  TL02_PHS1_knockback_mul_35_64_g1818 : MAOI22D0BWP7T port map(A1 => TL02_n_451, A2 => TL02_PHS1_knockback_mul_35_64_n_4, B1 => TL02_n_451, B2 => TL02_PHS1_knockback_mul_35_64_n_4, ZN => TL02_PHS1_knockback_mul_35_64_n_17);
  TL02_PHS1_knockback_mul_35_64_g1819 : MOAI22D0BWP7T port map(A1 => TL02_n_452, A2 => TL02_PHS1_knockback_mul_35_64_n_1, B1 => TL02_n_452, B2 => TL02_PHS1_knockback_mul_35_64_n_1, ZN => TL02_PHS1_knockback_mul_35_64_n_16);
  TL02_PHS1_knockback_mul_35_64_g1820 : MAOI22D0BWP7T port map(A1 => TL02_n_449, A2 => TL02_PHS1_knockback_mul_35_64_n_4, B1 => TL02_n_449, B2 => TL02_PHS1_knockback_mul_35_64_n_4, ZN => TL02_PHS1_knockback_mul_35_64_n_15);
  TL02_PHS1_knockback_mul_35_64_g1821 : MAOI22D0BWP7T port map(A1 => TL02_n_452, A2 => TL02_PHS1_knockback_mul_35_64_n_4, B1 => TL02_n_452, B2 => TL02_PHS1_knockback_mul_35_64_n_4, ZN => TL02_PHS1_knockback_mul_35_64_n_14);
  TL02_PHS1_knockback_mul_35_64_g1822 : MOAI22D0BWP7T port map(A1 => TL02_n_450, A2 => TL02_PHS1_knockback_mul_35_64_n_2, B1 => TL02_n_450, B2 => TL02_PHS1_knockback_mul_35_64_n_2, ZN => TL02_PHS1_knockback_mul_35_64_n_13);
  TL02_PHS1_knockback_mul_35_64_g1823 : MAOI22D0BWP7T port map(A1 => TL02_n_448, A2 => TL02_PHS1_knockback_mul_35_64_n_2, B1 => TL02_n_448, B2 => TL02_PHS1_knockback_mul_35_64_n_2, ZN => TL02_PHS1_knockback_mul_35_64_n_12);
  TL02_PHS1_knockback_mul_35_64_g1824 : MAOI22D0BWP7T port map(A1 => TL02_n_447, A2 => TL02_PHS1_knockback_mul_35_64_n_2, B1 => TL02_n_447, B2 => TL02_PHS1_knockback_mul_35_64_n_2, ZN => TL02_PHS1_knockback_mul_35_64_n_11);
  TL02_PHS1_knockback_mul_35_64_g1825 : MAOI22D0BWP7T port map(A1 => TL02_n_449, A2 => TL02_PHS1_knockback_mul_35_64_n_2, B1 => TL02_n_449, B2 => TL02_PHS1_knockback_mul_35_64_n_2, ZN => TL02_PHS1_knockback_mul_35_64_n_10);
  TL02_PHS1_knockback_mul_35_64_g1826 : MAOI22D0BWP7T port map(A1 => TL02_n_451, A2 => TL02_PHS1_knockback_mul_35_64_n_2, B1 => TL02_n_451, B2 => TL02_PHS1_knockback_mul_35_64_n_2, ZN => TL02_PHS1_knockback_mul_35_64_n_9);
  TL02_PHS1_knockback_mul_35_64_g1827 : MOAI22D0BWP7T port map(A1 => TL02_n_446, A2 => TL02_PHS1_knockback_mul_35_64_n_2, B1 => TL02_n_446, B2 => TL02_PHS1_knockback_mul_35_64_n_2, ZN => TL02_PHS1_knockback_mul_35_64_n_8);
  TL02_PHS1_knockback_mul_35_64_g1828 : INVD0BWP7T port map(I => TL02_PHS1_knockback_mul_35_64_n_7, ZN => TL02_PHS1_knockback_mul_35_64_n_6);
  TL02_PHS1_knockback_mul_35_64_g1829 : CKND2D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_5, A2 => TL02_n_444, ZN => TL02_PHS1_knockback_mul_35_64_n_7);
  TL02_PHS1_knockback_mul_35_64_g1830 : INVD1BWP7T port map(I => TL02_n_445, ZN => TL02_PHS1_knockback_mul_35_64_n_5);
  TL02_PHS1_knockback_mul_35_64_g1831 : INVD1BWP7T port map(I => TL02_n_438, ZN => TL02_PHS1_knockback_mul_35_64_n_4);
  TL02_PHS1_knockback_mul_35_64_g1832 : INVD1BWP7T port map(I => TL02_n_440, ZN => TL02_PHS1_knockback_mul_35_64_n_3);
  TL02_PHS1_knockback_mul_35_64_g1833 : INVD1BWP7T port map(I => TL02_n_444, ZN => TL02_PHS1_knockback_mul_35_64_n_2);
  TL02_PHS1_knockback_mul_35_64_g1834 : INVD1BWP7T port map(I => TL02_n_442, ZN => TL02_PHS1_knockback_mul_35_64_n_1);
  TL02_PHS1_knockback_mul_35_64_g1835 : XOR3D1BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_114, A2 => TL02_PHS1_knockback_mul_35_64_n_77, A3 => TL02_PHS1_knockback_mul_35_64_n_60, Z => TL02_PHS1_knockback_mul_35_64_n_199);
  TL02_PHS1_knockback_mul_35_64_g2 : OA21D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_106, A2 => TL02_PHS1_knockback_mul_35_64_n_200, B => TL02_PHS1_knockback_mul_35_64_n_57, Z => TL02_PHS1_knockback_mul_35_64_n_201);
  TL02_PHS1_knockback_mul_35_64_g3 : NR3D0BWP7T port map(A1 => TL02_PHS1_knockback_mul_35_64_n_2, A2 => TL02_n_453, A3 => TL02_n_452, ZN => TL02_PHS1_knockback_mul_35_64_n_200);
  TL01_g188 : INVD5BWP7T port map(I => TL01_n_63, ZN => Vsync);
  TL01_SCNR1_gen1_vgen_sync_reg : DFKSND1BWP7T port map(CP => CTS_17, D => FE_OFN3_reset, Q => UNCONNECTED, QN => TL01_n_63, SN => TL01_n_62);
  TL01_g191 : NR4D0BWP7T port map(A1 => TL01_n_59, A2 => vcountintern(2), A3 => vcountintern(1), A4 => vcountintern(9), ZN => TL01_n_62);
  TL01_g192 : AO21D0BWP7T port map(A1 => TL01_n_58, A2 => vcountintern(9), B => FE_OFN3_reset, Z => TL01_n_61);
  TL01_SCNR1_gen2_hgen_sync_reg : DFD1BWP7T port map(CP => CTS_16, D => TL01_n_57, Q => UNCONNECTED0, QN => TL01_n_60);
  TL01_g194 : INVD5BWP7T port map(I => TL01_n_60, ZN => Hsync);
  TL01_g195 : IND2D1BWP7T port map(A1 => vcountintern(3), B1 => TL01_n_56, ZN => TL01_n_59);
  TL01_g196 : ND2D1BWP7T port map(A1 => TL01_n_56, A2 => TL01_n_55, ZN => TL01_n_58);
  TL01_g197 : OR4D1BWP7T port map(A1 => FE_OFN3_reset, A2 => hcountintern(8), A3 => hcountintern(7), A4 => TL01_n_54, Z => TL01_n_57);
  TL01_g198 : NR4D0BWP7T port map(A1 => TL01_n_53, A2 => vcountintern(5), A3 => vcountintern(8), A4 => vcountintern(6), ZN => TL01_n_56);
  TL01_g199 : OAI211D1BWP7T port map(A1 => vcountintern(0), A2 => vcountintern(1), B => vcountintern(2), C => vcountintern(3), ZN => TL01_n_55);
  TL01_g200 : AO21D0BWP7T port map(A1 => hcountintern(5), A2 => hcountintern(6), B => hcountintern(9), Z => TL01_n_54);
  TL01_g201 : OR2D1BWP7T port map(A1 => vcountintern(4), A2 => vcountintern(7), Z => TL01_n_53);
  TL01_SCNR1_cnt1_vcnt_cur_count_reg_9 : DFKCNQD1BWP7T port map(CN => TL01_n_2, CP => CTS_16, D => TL01_n_52, Q => FE_PHN122_vcountintern_9);
  TL01_SCNR1_cnt1_vcnt_cur_count_reg_8 : DFKCNQD1BWP7T port map(CN => TL01_n_2, CP => CTS_16, D => TL01_n_50, Q => vcountintern(8));
  TL01_g370 : MOAI22D0BWP7T port map(A1 => TL01_n_49, A2 => TL01_n_15, B1 => TL01_n_15, B2 => vcountintern(9), ZN => TL01_n_52);
  TL01_g372 : MOAI22D0BWP7T port map(A1 => TL01_n_45, A2 => hcountintern(9), B1 => TL01_n_45, B2 => hcountintern(9), ZN => TL01_n_51);
  TL01_SCNR1_cnt2_hcnt_cur_count_reg_8 : DFKCNQD1BWP7T port map(CN => FE_PHN68_TL01_SCNR1_hcount_reset, CP => CTS_16, D => TL01_n_48, Q => hcountintern(8));
  TL01_g374 : MOAI22D0BWP7T port map(A1 => TL01_n_46, A2 => TL01_n_15, B1 => TL01_n_15, B2 => vcountintern(8), ZN => TL01_n_50);
  TL01_g375 : MAOI22D0BWP7T port map(A1 => TL01_n_44, A2 => vcountintern(9), B1 => TL01_n_44, B2 => vcountintern(9), ZN => TL01_n_49);
  TL01_SCNR1_cnt1_vcnt_cur_count_reg_7 : DFKCNQD1BWP7T port map(CN => TL01_n_2, CP => CTS_16, D => TL01_n_47, Q => vcountintern(7));
  TL01_g377 : MOAI22D0BWP7T port map(A1 => TL01_n_39, A2 => hcountintern(8), B1 => TL01_n_39, B2 => hcountintern(8), ZN => TL01_n_48);
  TL01_SCNR1_cnt2_hcnt_cur_count_reg_7 : DFKCNQD1BWP7T port map(CN => FE_PHN68_TL01_SCNR1_hcount_reset, CP => CTS_16, D => TL01_n_43, Q => hcountintern(7));
  TL01_g379 : MOAI22D0BWP7T port map(A1 => TL01_n_41, A2 => TL01_n_15, B1 => TL01_n_15, B2 => vcountintern(7), ZN => TL01_n_47);
  TL01_g380 : MAOI22D0BWP7T port map(A1 => TL01_n_40, A2 => vcountintern(8), B1 => TL01_n_40, B2 => vcountintern(8), ZN => TL01_n_46);
  TL01_SCNR1_cnt1_vcnt_cur_count_reg_6 : DFKCNQD1BWP7T port map(CN => TL01_n_2, CP => CTS_16, D => TL01_n_42, Q => vcountintern(6));
  TL01_g382 : IND2D1BWP7T port map(A1 => TL01_n_39, B1 => hcountintern(8), ZN => TL01_n_45);
  TL01_g383 : IND2D1BWP7T port map(A1 => TL01_n_40, B1 => vcountintern(8), ZN => TL01_n_44);
  TL01_g384 : MOAI22D0BWP7T port map(A1 => TL01_n_34, A2 => hcountintern(7), B1 => TL01_n_34, B2 => hcountintern(7), ZN => TL01_n_43);
  TL01_SCNR1_cnt2_hcnt_cur_count_reg_6 : DFKCNQD1BWP7T port map(CN => FE_PHN68_TL01_SCNR1_hcount_reset, CP => CTS_16, D => TL01_n_38, Q => hcountintern(6));
  TL01_g386 : MOAI22D0BWP7T port map(A1 => TL01_n_36, A2 => TL01_n_15, B1 => TL01_n_15, B2 => vcountintern(6), ZN => TL01_n_42);
  TL01_g387 : MAOI22D0BWP7T port map(A1 => TL01_n_35, A2 => vcountintern(7), B1 => TL01_n_35, B2 => vcountintern(7), ZN => TL01_n_41);
  TL01_SCNR1_cnt1_vcnt_cur_count_reg_5 : DFKCNQD1BWP7T port map(CN => TL01_n_2, CP => CTS_16, D => TL01_n_37, Q => vcountintern(5));
  TL01_g389 : IND2D1BWP7T port map(A1 => TL01_n_35, B1 => vcountintern(7), ZN => TL01_n_40);
  TL01_g390 : IND2D1BWP7T port map(A1 => TL01_n_34, B1 => hcountintern(7), ZN => TL01_n_39);
  TL01_g391 : MOAI22D0BWP7T port map(A1 => TL01_n_30, A2 => hcountintern(6), B1 => TL01_n_30, B2 => hcountintern(6), ZN => TL01_n_38);
  TL01_SCNR1_cnt2_hcnt_cur_count_reg_5 : DFKCNQD1BWP7T port map(CN => FE_PHN68_TL01_SCNR1_hcount_reset, CP => CTS_16, D => TL01_n_32, Q => hcountintern(5));
  TL01_g393 : MOAI22D0BWP7T port map(A1 => TL01_n_15, A2 => TL01_n_31, B1 => TL01_n_15, B2 => vcountintern(5), ZN => TL01_n_37);
  TL01_g394 : MAOI22D0BWP7T port map(A1 => TL01_n_29, A2 => vcountintern(6), B1 => TL01_n_29, B2 => vcountintern(6), ZN => TL01_n_36);
  TL01_SCNR1_cnt1_vcnt_cur_count_reg_4 : DFKCNQD1BWP7T port map(CN => TL01_n_2, CP => CTS_16, D => TL01_n_33, Q => vcountintern(4));
  TL01_g396 : IND2D1BWP7T port map(A1 => TL01_n_29, B1 => vcountintern(6), ZN => TL01_n_35);
  TL01_g397 : IND2D1BWP7T port map(A1 => TL01_n_30, B1 => hcountintern(6), ZN => TL01_n_34);
  TL01_g398 : MOAI22D0BWP7T port map(A1 => TL01_n_15, A2 => TL01_n_28, B1 => TL01_n_15, B2 => vcountintern(4), ZN => TL01_n_33);
  TL01_SCNR1_cnt2_hcnt_cur_count_reg_4 : DFKCNQD1BWP7T port map(CN => FE_PHN68_TL01_SCNR1_hcount_reset, CP => CTS_16, D => TL01_n_27, Q => hcountintern(4));
  TL01_g400 : MOAI22D0BWP7T port map(A1 => TL01_n_25, A2 => hcountintern(5), B1 => TL01_n_25, B2 => hcountintern(5), ZN => TL01_n_32);
  TL01_g401 : MAOI22D0BWP7T port map(A1 => TL01_n_24, A2 => vcountintern(5), B1 => TL01_n_24, B2 => vcountintern(5), ZN => TL01_n_31);
  TL01_SCNR1_cnt1_vcnt_cur_count_reg_3 : DFKCNQD1BWP7T port map(CN => TL01_n_2, CP => CTS_16, D => TL01_n_26, Q => vcountintern(3));
  TL01_g403 : IND2D1BWP7T port map(A1 => TL01_n_25, B1 => hcountintern(5), ZN => TL01_n_30);
  TL01_g404 : IND2D1BWP7T port map(A1 => TL01_n_24, B1 => vcountintern(5), ZN => TL01_n_29);
  TL01_SCNR1_cnt1_vcnt_cur_count_reg_1 : DFKCNQD1BWP7T port map(CN => TL01_n_2, CP => CTS_16, D => TL01_n_23, Q => vcountintern(1));
  TL01_SCNR1_cnt1_vcnt_cur_count_reg_2 : DFKCNQD1BWP7T port map(CN => TL01_n_2, CP => CTS_16, D => TL01_n_21, Q => vcountintern(2));
  TL01_SCNR1_cnt1_vcnt_cur_count_reg_0 : DFKCNQD1BWP7T port map(CN => TL01_n_2, CP => CTS_16, D => TL01_n_22, Q => vcountintern(0));
  TL01_g408 : MAOI22D0BWP7T port map(A1 => TL01_n_16, A2 => vcountintern(4), B1 => TL01_n_16, B2 => vcountintern(4), ZN => TL01_n_28);
  TL01_g409 : MOAI22D0BWP7T port map(A1 => TL01_n_17, A2 => hcountintern(4), B1 => TL01_n_17, B2 => hcountintern(4), ZN => TL01_n_27);
  TL01_g410 : MOAI22D0BWP7T port map(A1 => TL01_n_15, A2 => TL01_n_18, B1 => TL01_n_15, B2 => vcountintern(3), ZN => TL01_n_26);
  TL01_SCNR1_cnt2_hcnt_cur_count_reg_3 : DFKCNQD1BWP7T port map(CN => FE_PHN68_TL01_SCNR1_hcount_reset, CP => CTS_16, D => TL01_n_19, Q => hcountintern(3));
  TL01_g412 : IND2D1BWP7T port map(A1 => TL01_n_17, B1 => hcountintern(4), ZN => TL01_n_25);
  TL01_g413 : IND2D1BWP7T port map(A1 => TL01_n_16, B1 => vcountintern(4), ZN => TL01_n_24);
  TL01_g414 : MOAI22D0BWP7T port map(A1 => TL01_n_15, A2 => TL01_n_6, B1 => TL01_n_15, B2 => vcountintern(1), ZN => TL01_n_23);
  TL01_SCNR1_gen2_hgen_cnt_reset_reg : DFD1BWP7T port map(CP => CTS_16, D => TL01_n_20, Q => UNCONNECTED1, QN => TL01_SCNR1_hcount_reset);
  TL01_g416 : MOAI22D0BWP7T port map(A1 => TL01_n_15, A2 => vcountintern(0), B1 => TL01_n_15, B2 => vcountintern(0), ZN => TL01_n_22);
  TL01_g417 : MOAI22D0BWP7T port map(A1 => TL01_n_15, A2 => TL01_n_12, B1 => TL01_n_15, B2 => vcountintern(2), ZN => TL01_n_21);
  TL01_g418 : AO211D0BWP7T port map(A1 => TL01_n_11, A2 => hcountintern(8), B => TL01_n_14, C => FE_OFN3_reset, Z => TL01_n_20);
  TL01_SCNR1_cnt2_hcnt_cur_count_reg_2 : DFKCNQD1BWP7T port map(CN => FE_PHN68_TL01_SCNR1_hcount_reset, CP => CTS_16, D => TL01_n_13, Q => hcountintern(2));
  TL01_g420 : MOAI22D0BWP7T port map(A1 => TL01_n_9, A2 => hcountintern(3), B1 => TL01_n_9, B2 => hcountintern(3), ZN => TL01_n_19);
  TL01_g421 : MAOI22D0BWP7T port map(A1 => TL01_n_10, A2 => vcountintern(3), B1 => TL01_n_10, B2 => vcountintern(3), ZN => TL01_n_18);
  TL01_g422 : IND2D1BWP7T port map(A1 => TL01_n_9, B1 => hcountintern(3), ZN => TL01_n_17);
  TL01_g423 : IND2D1BWP7T port map(A1 => TL01_n_10, B1 => vcountintern(3), ZN => TL01_n_16);
  TL01_g424 : IND3D1BWP7T port map(A1 => TL01_hcount_int(0), B1 => TL01_n_7, B2 => TL01_n_14, ZN => TL01_n_15);
  TL01_g425 : AN3D1BWP7T port map(A1 => TL01_n_8, A2 => hcountintern(1), A3 => hcountintern(8), Z => TL01_n_14);
  TL01_SCNR1_cnt2_hcnt_cur_count_reg_1 : DFKCNQD1BWP7T port map(CN => FE_PHN68_TL01_SCNR1_hcount_reset, CP => CTS_16, D => TL01_n_5, Q => hcountintern(1));
  TL01_g427 : MOAI22D0BWP7T port map(A1 => TL01_n_4, A2 => hcountintern(2), B1 => TL01_n_4, B2 => hcountintern(2), ZN => TL01_n_13);
  TL01_g428 : MAOI22D0BWP7T port map(A1 => TL01_n_3, A2 => vcountintern(2), B1 => TL01_n_3, B2 => vcountintern(2), ZN => TL01_n_12);
  TL01_g429 : MOAI22D0BWP7T port map(A1 => TL01_n_7, A2 => FE_PHN96_TL01_n_1, B1 => TL01_n_8, B2 => TL01_hcount_int(0), ZN => TL01_n_11);
  TL01_g430 : IND2D1BWP7T port map(A1 => TL01_n_3, B1 => vcountintern(2), ZN => TL01_n_10);
  TL01_g431 : IND2D1BWP7T port map(A1 => TL01_n_4, B1 => hcountintern(2), ZN => TL01_n_9);
  TL01_g432 : AN4D1BWP7T port map(A1 => hcountintern(3), A2 => hcountintern(2), A3 => hcountintern(9), A4 => hcountintern(4), Z => TL01_n_8);
  TL01_g433 : NR3D0BWP7T port map(A1 => hcountintern(5), A2 => hcountintern(6), A3 => hcountintern(7), ZN => TL01_n_7);
  TL01_g435 : XNR2D1BWP7T port map(A1 => vcountintern(0), A2 => vcountintern(1), ZN => TL01_n_6);
  TL01_g436 : MOAI22D0BWP7T port map(A1 => TL01_n_0, A2 => hcountintern(1), B1 => TL01_n_0, B2 => hcountintern(1), ZN => TL01_n_5);
  TL01_g437 : ND2D1BWP7T port map(A1 => TL01_hcount_int(0), A2 => hcountintern(1), ZN => TL01_n_4);
  TL01_g438 : ND2D1BWP7T port map(A1 => vcountintern(1), A2 => vcountintern(0), ZN => TL01_n_3);
  TL01_SCNR1_gen1_vgen_cnt_reset_reg : DFD1BWP7T port map(CP => CTS_16, D => TL01_n_61, Q => TL01_SCNR1_vcount_reset, QN => FE_PHN34_TL01_n_2);
  TL01_SCNR1_cnt2_hcnt_cur_count_reg_9 : DFKCND1BWP7T port map(CN => FE_PHN68_TL01_SCNR1_hcount_reset, CP => CTS_16, D => TL01_n_51, Q => hcountintern(9), QN => TL01_n_1);
  TL01_SCNR1_cnt2_hcnt_cur_count_reg_0 : DFKCND1BWP7T port map(CN => FE_PHN158_TL01_n_0, CP => CTS_16, D => FE_PHN160_TL01_SCNR1_hcount_reset, Q => TL01_hcount_int(0), QN => FE_PHN62_TL01_n_0);
  TL01_CLR1_B_data_reg_0 : DFD0BWP7T port map(CP => CTS_16, D => TL01_CLR1_n_1456, Q => UNCONNECTED2, QN => TL01_CLR1_n_1464);
  TL01_CLR1_B_data_reg_1 : DFD0BWP7T port map(CP => CTS_16, D => TL01_CLR1_n_1454, Q => UNCONNECTED3, QN => TL01_CLR1_n_1461);
  TL01_CLR1_B_data_reg_2 : DFD0BWP7T port map(CP => CTS_16, D => TL01_CLR1_n_1469, Q => UNCONNECTED4, QN => TL01_CLR1_n_1473);
  TL01_CLR1_B_data_reg_3 : DFD0BWP7T port map(CP => CTS_16, D => TL01_CLR1_n_1468, Q => UNCONNECTED5, QN => TL01_CLR1_n_1470);
  TL01_CLR1_G_data_reg_0 : DFD0BWP7T port map(CP => CTS_16, D => TL01_CLR1_n_1467, Q => UNCONNECTED6, QN => TL01_CLR1_n_1471);
  TL01_CLR1_G_data_reg_1 : DFD0BWP7T port map(CP => CTS_16, D => TL01_CLR1_n_1457, Q => UNCONNECTED7, QN => TL01_CLR1_n_1460);
  TL01_CLR1_G_data_reg_2 : DFD0BWP7T port map(CP => CTS_16, D => TL01_CLR1_n_1452, Q => UNCONNECTED8, QN => TL01_CLR1_n_1459);
  TL01_CLR1_R_data_reg_0 : DFD0BWP7T port map(CP => CTS_16, D => TL01_CLR1_n_1455, Q => UNCONNECTED9, QN => TL01_CLR1_n_1463);
  TL01_CLR1_R_data_reg_2 : DFD0BWP7T port map(CP => CTS_16, D => TL01_CLR1_n_1466, Q => UNCONNECTED10, QN => TL01_CLR1_n_1472);
  TL01_CLR1_char1_sprite_frame_control_new_state_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => FE_PHN144_TL01_CLR1_n_733, Q => TL01_CLR1_char1_sprite_frame_control_new_state_0);
  TL01_CLR1_char1_sprite_frame_control_new_state_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL01_CLR1_n_672, Q => TL01_CLR1_char1_sprite_frame_control_new_state_1);
  TL01_CLR1_char1_sprite_frame_control_new_state_reg_2 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL01_CLR1_n_704, Q => TL01_CLR1_char1_sprite_frame_control_new_state_2);
  TL01_CLR1_char1_sprite_frame_control_sprite_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL01_CLR1_n_3, Q => TL01_CLR1_char1_sprite_sprite_1);
  TL01_CLR1_char2_sprite_frame_control_new_state_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_15, D => TL01_CLR1_n_737, Q => TL01_CLR1_char2_sprite_frame_control_new_state_0);
  TL01_CLR1_char2_sprite_frame_control_new_state_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_15, D => TL01_CLR1_n_671, Q => TL01_CLR1_char2_sprite_frame_control_new_state_1);
  TL01_CLR1_char2_sprite_frame_control_new_state_reg_2 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_15, D => TL01_CLR1_n_703, Q => TL01_CLR1_char2_sprite_frame_control_new_state_2);
  TL01_CLR1_char2_sprite_frame_control_sprite_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => FE_PHN152_TL01_CLR1_n_303, Q => TL01_CLR1_char2_sprite_sprite_0);
  TL01_CLR1_char2_sprite_frame_control_sprite_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL01_CLR1_n_2, Q => TL01_CLR1_char2_sprite_sprite_1);
  TL01_CLR1_g40524 : CKND10BWP7T port map(I => TL01_CLR1_n_1473, ZN => G_data(3));
  TL01_CLR1_g40526 : CKND10BWP7T port map(I => TL01_CLR1_n_1472, ZN => R_data(3));
  TL01_CLR1_g40528 : INVD5BWP7T port map(I => TL01_CLR1_n_1471, ZN => G_data(0));
  TL01_CLR1_g40530 : INVD5BWP7T port map(I => TL01_CLR1_n_1470, ZN => B_data(3));
  TL01_CLR1_g40531 : IND4D0BWP7T port map(A1 => TL01_CLR1_n_1450, B1 => TL01_CLR1_n_1444, B2 => TL01_CLR1_n_1435, B3 => TL01_CLR1_n_1465, ZN => TL01_CLR1_n_1469);
  TL01_CLR1_g40532 : IND4D0BWP7T port map(A1 => TL01_CLR1_n_1450, B1 => TL01_CLR1_n_1425, B2 => TL01_CLR1_n_1443, B3 => TL01_CLR1_n_1465, ZN => TL01_CLR1_n_1468);
  TL01_CLR1_g40533 : ND4D0BWP7T port map(A1 => TL01_CLR1_n_1462, A2 => TL01_CLR1_n_1442, A3 => TL01_CLR1_n_1246, A4 => TL01_CLR1_n_1449, ZN => TL01_CLR1_n_1467);
  TL01_CLR1_g40534 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_1465, A2 => TL01_CLR1_n_1246, A3 => TL01_CLR1_n_1449, ZN => TL01_CLR1_n_1466);
  TL01_CLR1_g40535 : INR2XD0BWP7T port map(A1 => TL01_CLR1_n_1462, B1 => TL01_CLR1_n_1446, ZN => TL01_CLR1_n_1465);
  TL01_CLR1_g40537 : INVD5BWP7T port map(I => TL01_CLR1_n_1464, ZN => B_data(0));
  TL01_CLR1_g40539 : INVD5BWP7T port map(I => TL01_CLR1_n_1463, ZN => R_data(0));
  TL01_CLR1_g40541 : INVD5BWP7T port map(I => TL01_CLR1_n_1461, ZN => B_data(1));
  TL01_CLR1_g40543 : CKND10BWP7T port map(I => TL01_CLR1_n_1460, ZN => R_data(1));
  TL01_CLR1_g40544 : AOI211XD0BWP7T port map(A1 => TL01_CLR1_n_1448, A2 => hcountintern(7), B => TL01_CLR1_n_1458, C => TL01_CLR1_n_1447, ZN => TL01_CLR1_n_1462);
  TL01_CLR1_g40546 : INVD5BWP7T port map(I => TL01_CLR1_n_1459, ZN => G_data(2));
  TL01_CLR1_g40547 : OAI31D0BWP7T port map(A1 => hcountintern(9), A2 => TL01_CLR1_n_154, A3 => TL01_CLR1_n_1436, B => TL01_CLR1_n_1453, ZN => TL01_CLR1_n_1458);
  TL01_CLR1_g40548 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_1451, A2 => TL01_CLR1_n_1246, A3 => TL01_CLR1_n_1444, ZN => TL01_CLR1_n_1457);
  TL01_CLR1_g40549 : IND4D0BWP7T port map(A1 => TL01_CLR1_n_1450, B1 => TL01_CLR1_n_1449, B2 => TL01_CLR1_n_1438, B3 => TL01_CLR1_n_1442, ZN => TL01_CLR1_n_1456);
  TL01_CLR1_g40550 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_1442, A2 => TL01_CLR1_n_49, A3 => TL01_CLR1_n_1444, ZN => TL01_CLR1_n_1455);
  TL01_CLR1_g40551 : IND3D1BWP7T port map(A1 => TL01_CLR1_n_1450, B1 => TL01_CLR1_n_1444, B2 => TL01_CLR1_n_1451, ZN => TL01_CLR1_n_1454);
  TL01_CLR1_g40552 : AOI32D1BWP7T port map(A1 => TL01_CLR1_n_1437, A2 => TL01_CLR1_n_157, A3 => hcountintern(9), B1 => TL01_CLR1_n_1439, B2 => TL01_CLR1_n_691, ZN => TL01_CLR1_n_1453);
  TL01_CLR1_g40553 : IND3D1BWP7T port map(A1 => TL01_CLR1_n_1445, B1 => TL01_CLR1_n_1444, B2 => TL01_CLR1_n_1440, ZN => TL01_CLR1_n_1452);
  TL01_CLR1_g40555 : INR2XD0BWP7T port map(A1 => TL01_CLR1_n_1438, B1 => TL01_CLR1_n_1446, ZN => TL01_CLR1_n_1451);
  TL01_CLR1_g40556 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1246, A2 => TL01_CLR1_n_1441, ZN => TL01_CLR1_n_1450);
  TL01_CLR1_g40557 : NR4D0BWP7T port map(A1 => TL01_CLR1_n_1403, A2 => TL01_CLR1_n_1430, A3 => TL01_CLR1_n_81, A4 => hcountintern(6), ZN => TL01_CLR1_n_1448);
  TL01_CLR1_g40558 : AN4D0BWP7T port map(A1 => TL01_CLR1_n_1427, A2 => TL01_CLR1_n_1424, A3 => TL01_CLR1_n_837, A4 => TL01_CLR1_n_364, Z => TL01_CLR1_n_1447);
  TL01_CLR1_g40559 : OA21D0BWP7T port map(A1 => TL01_CLR1_n_1417, A2 => TL01_CLR1_n_1364, B => TL01_CLR1_n_1443, Z => TL01_CLR1_n_1449);
  TL01_CLR1_g40560 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1440, A2 => TL01_CLR1_n_1433, ZN => TL01_CLR1_n_1446);
  TL01_CLR1_g40561 : INR4D0BWP7T port map(A1 => TL01_CLR1_n_1417, B1 => TL01_CLR1_n_1431, B2 => TL01_CLR1_n_916, B3 => TL01_CLR1_n_1428, ZN => TL01_CLR1_n_1445);
  TL01_CLR1_g40562 : OA21D0BWP7T port map(A1 => TL01_CLR1_n_1432, A2 => TL01_CLR1_n_1341, B => TL01_CLR1_n_1425, Z => TL01_CLR1_n_1444);
  TL01_CLR1_g40563 : AOI211XD0BWP7T port map(A1 => TL01_CLR1_n_1424, A2 => TL01_CLR1_n_692, B => TL01_CLR1_n_1429, C => TL01_CLR1_n_1418, ZN => TL01_CLR1_n_1441);
  TL01_CLR1_g40564 : OA21D0BWP7T port map(A1 => TL01_CLR1_n_1432, A2 => TL01_CLR1_n_1226, B => TL01_CLR1_n_1435, Z => TL01_CLR1_n_1443);
  TL01_CLR1_g40565 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1428, A2 => TL01_CLR1_n_768, B1 => TL01_CLR1_n_1434, B2 => TL01_CLR1_n_514, ZN => TL01_CLR1_n_1442);
  TL01_CLR1_g40566 : AOI211D1BWP7T port map(A1 => TL01_CLR1_n_1419, A2 => TL01_CLR1_n_1281, B => TL01_CLR1_n_1422, C => TL01_CLR1_n_439, ZN => TL01_CLR1_n_1439);
  TL01_CLR1_g40567 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1428, A2 => TL01_CLR1_n_1351, ZN => TL01_CLR1_n_1440);
  TL01_CLR1_g40568 : AOI211D1BWP7T port map(A1 => TL01_CLR1_n_1493, A2 => TL01_CLR1_n_146, B => TL01_CLR1_n_1412, C => TL01_CLR1_n_1430, ZN => TL01_CLR1_n_1437);
  TL01_CLR1_g40569 : AO211D0BWP7T port map(A1 => TL01_CLR1_n_496, A2 => TL01_CLR1_n_1493, B => TL01_CLR1_n_1415, C => TL01_CLR1_n_1430, Z => TL01_CLR1_n_1436);
  TL01_CLR1_g40570 : OA21D0BWP7T port map(A1 => TL01_CLR1_n_1423, A2 => TL01_CLR1_n_1332, B => TL01_CLR1_n_1422, Z => TL01_CLR1_n_1438);
  TL01_CLR1_g40571 : INVD0BWP7T port map(I => TL01_CLR1_n_1433, ZN => TL01_CLR1_n_1434);
  TL01_CLR1_g40572 : CKND1BWP7T port map(I => TL01_CLR1_n_1431, ZN => TL01_CLR1_n_1432);
  TL01_CLR1_g40573 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_1405, A2 => TL01_CLR1_n_1424, A3 => TL01_CLR1_n_837, ZN => TL01_CLR1_n_1435);
  TL01_CLR1_g40574 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1424, A2 => TL01_CLR1_n_1270, ZN => TL01_CLR1_n_1433);
  TL01_CLR1_g40575 : NR3D0BWP7T port map(A1 => TL01_CLR1_n_1420, A2 => TL01_CLR1_n_1413, A3 => TL01_CLR1_n_47, ZN => TL01_CLR1_n_1431);
  TL01_CLR1_g40576 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1424, A2 => TL01_CLR1_n_691, ZN => TL01_CLR1_n_1430);
  TL01_CLR1_g40578 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_1179, A2 => TL01_CLR1_n_1037, B1 => TL01_CLR1_n_1036, B2 => TL01_CLR1_n_1120, C => TL01_CLR1_n_1421, ZN => TL01_CLR1_n_1427);
  TL01_CLR1_g40579 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_1270, A2 => TL01_CLR1_n_692, B => TL01_CLR1_n_1424, ZN => TL01_CLR1_n_1426);
  TL01_CLR1_g40580 : INR3D0BWP7T port map(A1 => TL01_CLR1_n_47, B1 => TL01_CLR1_n_1413, B2 => TL01_CLR1_n_1420, ZN => TL01_CLR1_n_1429);
  TL01_CLR1_g40581 : NR3D0BWP7T port map(A1 => TL01_CLR1_n_1423, A2 => TL01_CLR1_n_1306, A3 => TL01_CLR1_n_806, ZN => TL01_CLR1_n_1428);
  TL01_CLR1_g40582 : INVD0BWP7T port map(I => TL01_CLR1_n_1424, ZN => TL01_CLR1_n_1423);
  TL01_CLR1_g40583 : IND4D0BWP7T port map(A1 => TL01_CLR1_n_1417, B1 => TL01_CLR1_n_575, B2 => TL01_CLR1_n_1257, B3 => TL01_CLR1_n_1018, ZN => TL01_CLR1_n_1425);
  TL01_CLR1_g40584 : INR2XD0BWP7T port map(A1 => TL01_CLR1_n_1413, B1 => TL01_CLR1_n_1420, ZN => TL01_CLR1_n_1424);
  TL01_CLR1_g40585 : AOI31D0BWP7T port map(A1 => TL01_CLR1_n_1089, A2 => TL01_CLR1_n_1034, A3 => TL01_CLR1_n_310, B => TL01_CLR1_n_1416, ZN => TL01_CLR1_n_1421);
  TL01_CLR1_g40586 : IND3D1BWP7T port map(A1 => TL01_CLR1_n_1137, B1 => TL01_CLR1_n_1413, B2 => TL01_CLR1_n_1414, ZN => TL01_CLR1_n_1422);
  TL01_CLR1_g40587 : NR4D0BWP7T port map(A1 => TL01_CLR1_n_1409, A2 => TL01_CLR1_n_1389, A3 => TL01_CLR1_n_1284, A4 => TL01_CLR1_n_1202, ZN => TL01_CLR1_n_1419);
  TL01_CLR1_g40588 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1414, A2 => TL01_CLR1_n_1222, ZN => TL01_CLR1_n_1420);
  TL01_CLR1_g40589 : IND4D0BWP7T port map(A1 => TL01_CLR1_n_1384, B1 => TL01_CLR1_n_1176, B2 => TL01_CLR1_n_1309, B3 => TL01_CLR1_n_1411, ZN => TL01_CLR1_n_1416);
  TL01_CLR1_g40590 : INR3D0BWP7T port map(A1 => TL01_CLR1_n_1222, B1 => TL01_CLR1_n_1378, B2 => TL01_CLR1_n_1414, ZN => TL01_CLR1_n_1418);
  TL01_CLR1_g40591 : IND3D1BWP7T port map(A1 => TL01_CLR1_n_1414, B1 => TL01_CLR1_n_1378, B2 => TL01_CLR1_n_1222, ZN => TL01_CLR1_n_1417);
  TL01_CLR1_g40592 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_496, A2 => TL01_CLR1_n_124, B => TL01_CLR1_n_1410, ZN => TL01_CLR1_n_1415);
  TL01_CLR1_g40593 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_1365, A2 => TL01_CLR1_n_1369, B => TL01_CLR1_n_1408, C => TL01_CLR1_n_1404, ZN => TL01_CLR1_n_1414);
  TL01_CLR1_g40594 : OAI32D1BWP7T port map(A1 => TL01_CLR1_n_1344, A2 => TL01_CLR1_n_1390, A3 => TL01_CLR1_n_1401, B1 => TL01_CLR1_n_167, B2 => TL01_CLR1_n_146, ZN => TL01_CLR1_n_1412);
  TL01_CLR1_g40595 : ND4D0BWP7T port map(A1 => TL01_CLR1_n_1402, A2 => TL01_CLR1_n_1395, A3 => TL01_CLR1_n_1393, A4 => TL01_CLR1_n_1381, ZN => TL01_CLR1_n_1413);
  TL01_CLR1_g40596 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_1031, A2 => TL01_CLR1_n_854, B1 => TL01_CLR1_n_1068, B2 => TL01_CLR1_n_682, C => TL01_CLR1_n_1407, ZN => TL01_CLR1_n_1411);
  TL01_CLR1_g40597 : AO211D0BWP7T port map(A1 => TL01_CLR1_n_1174, A2 => TL01_CLR1_n_1102, B => TL01_CLR1_n_1406, C => TL01_CLR1_n_1391, Z => TL01_CLR1_n_1410);
  TL01_CLR1_g40598 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_908, A2 => TL01_CLR1_n_1153, B => TL01_CLR1_n_1399, C => TL01_CLR1_n_1297, ZN => TL01_CLR1_n_1409);
  TL01_CLR1_g40599 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1398, A2 => vcountintern(9), B1 => TL01_CLR1_n_1386, B2 => TL01_CLR1_n_1167, ZN => TL01_CLR1_n_1408);
  TL01_CLR1_g40600 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_993, A2 => TL01_CLR1_n_1030, B1 => TL01_CLR1_n_903, B2 => TL01_CLR1_n_1096, C => TL01_CLR1_n_1400, ZN => TL01_CLR1_n_1407);
  TL01_CLR1_g40601 : ND4D0BWP7T port map(A1 => TL01_CLR1_n_1396, A2 => TL01_CLR1_n_1376, A3 => TL01_CLR1_n_1283, A4 => TL01_CLR1_n_1237, ZN => TL01_CLR1_n_1406);
  TL01_CLR1_g40602 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_496, A2 => TL01_CLR1_n_168, B => TL01_CLR1_n_1397, ZN => TL01_CLR1_n_1405);
  TL01_CLR1_g40603 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_1379, A2 => TL01_CLR1_n_81, B1 => TL01_CLR1_n_1392, B2 => TL01_CLR1_n_1331, C1 => TL01_CLR1_n_1373, C2 => TL01_CLR1_n_1291, ZN => TL01_CLR1_n_1404);
  TL01_CLR1_g40604 : OAI222D0BWP7T port map(A1 => TL01_CLR1_n_1387, A2 => TL01_CLR1_n_1282, B1 => TL01_CLR1_n_124, B2 => TL01_CLR1_n_150, C1 => TL01_CLR1_n_101, C2 => TL01_CLR1_n_149, ZN => TL01_CLR1_n_1403);
  TL01_CLR1_g40605 : AOI31D0BWP7T port map(A1 => TL01_CLR1_n_1298, A2 => TL01_CLR1_n_1301, A3 => TL01_CLR1_n_1293, B => TL01_CLR1_n_1394, ZN => TL01_CLR1_n_1402);
  TL01_CLR1_g40606 : IND4D0BWP7T port map(A1 => TL01_CLR1_n_1371, B1 => TL01_CLR1_n_1296, B2 => TL01_CLR1_n_1352, B3 => TL01_CLR1_n_1368, ZN => TL01_CLR1_n_1401);
  TL01_CLR1_g40607 : AOI211XD0BWP7T port map(A1 => TL01_CLR1_n_1128, A2 => TL01_CLR1_n_489, B => TL01_CLR1_n_1388, C => TL01_CLR1_n_1380, ZN => TL01_CLR1_n_1400);
  TL01_CLR1_g40608 : NR4D0BWP7T port map(A1 => TL01_CLR1_n_1385, A2 => TL01_CLR1_n_1357, A3 => TL01_CLR1_n_1330, A4 => TL01_CLR1_n_1245, ZN => TL01_CLR1_n_1399);
  TL01_CLR1_g40609 : OA211D0BWP7T port map(A1 => TL01_CLR1_n_147, A2 => TL01_CLR1_n_1200, B => TL01_CLR1_n_1386, C => TL01_CLR1_n_1167, Z => TL01_CLR1_n_1398);
  TL01_CLR1_g40610 : OAI31D0BWP7T port map(A1 => TL01_CLR1_n_1265, A2 => TL01_CLR1_n_1367, A3 => TL01_CLR1_n_1374, B => TL01_CLR1_n_670, ZN => TL01_CLR1_n_1397);
  TL01_CLR1_g40611 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_1092, A2 => TL01_CLR1_n_856, B1 => TL01_CLR1_n_1098, B2 => TL01_CLR1_n_656, C => TL01_CLR1_n_1383, ZN => TL01_CLR1_n_1396);
  TL01_CLR1_g40612 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_1170, A2 => TL01_CLR1_n_147, B1 => vcountintern(9), B2 => TL01_CLR1_n_1163, C => TL01_CLR1_n_1382, ZN => TL01_CLR1_n_1395);
  TL01_CLR1_g40613 : OA21D0BWP7T port map(A1 => TL01_CLR1_n_1377, A2 => TL01_CLR1_n_81, B => TL01_CLR1_n_1333, Z => TL01_CLR1_n_1394);
  TL01_CLR1_g40614 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1377, A2 => TL01_CLR1_n_81, B1 => TL01_CLR1_n_1227, B2 => TL01_CLR1_n_148, ZN => TL01_CLR1_n_1393);
  TL01_CLR1_g40615 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_1379, A2 => TL01_CLR1_n_81, Z => TL01_CLR1_n_1392);
  TL01_CLR1_g40616 : ND4D0BWP7T port map(A1 => TL01_CLR1_n_1372, A2 => TL01_CLR1_n_1350, A3 => TL01_CLR1_n_1342, A4 => TL01_CLR1_n_1241, ZN => TL01_CLR1_n_1391);
  TL01_CLR1_g40617 : ND4D0BWP7T port map(A1 => TL01_CLR1_n_1359, A2 => TL01_CLR1_n_1343, A3 => TL01_CLR1_n_1340, A4 => TL01_CLR1_n_1276, ZN => TL01_CLR1_n_1390);
  TL01_CLR1_g40618 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_387, A2 => TL01_CLR1_n_1263, B => TL01_CLR1_n_1362, C => TL01_CLR1_n_1360, ZN => TL01_CLR1_n_1389);
  TL01_CLR1_g40619 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_892, A2 => TL01_CLR1_n_1096, B => TL01_CLR1_n_1366, C => TL01_CLR1_n_1313, ZN => TL01_CLR1_n_1388);
  TL01_CLR1_g40620 : IND4D0BWP7T port map(A1 => TL01_CLR1_n_1310, B1 => TL01_CLR1_n_893, B2 => TL01_CLR1_n_1125, B3 => TL01_CLR1_n_1375, ZN => TL01_CLR1_n_1387);
  TL01_CLR1_g40621 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_1088, A2 => TL01_CLR1_n_881, B1 => TL01_CLR1_n_1114, B2 => TL01_CLR1_n_1308, C => TL01_CLR1_n_1353, ZN => TL01_CLR1_n_1385);
  TL01_CLR1_g40622 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_1037, A2 => TL01_CLR1_n_989, B => TL01_CLR1_n_1355, C => TL01_CLR1_n_1290, ZN => TL01_CLR1_n_1384);
  TL01_CLR1_g40623 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_863, A2 => TL01_CLR1_n_1091, B => TL01_CLR1_n_1358, C => TL01_CLR1_n_1320, ZN => TL01_CLR1_n_1383);
  TL01_CLR1_g40624 : OAI31D0BWP7T port map(A1 => TL01_CLR1_n_1256, A2 => TL01_CLR1_n_1295, A3 => TL01_CLR1_n_1346, B => TL01_CLR1_n_1292, ZN => TL01_CLR1_n_1382);
  TL01_CLR1_g40625 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1323, A2 => TL01_CLR1_n_1354, B1 => TL01_CLR1_n_1363, B2 => TL01_CLR1_n_123, ZN => TL01_CLR1_n_1381);
  TL01_CLR1_g40626 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_236, A2 => TL01_CLR1_n_1212, B => TL01_CLR1_n_1361, C => TL01_CLR1_n_1255, ZN => TL01_CLR1_n_1380);
  TL01_CLR1_g40627 : IOA21D1BWP7T port map(A1 => TL01_CLR1_n_1200, A2 => vcountintern(8), B => TL01_CLR1_n_1370, ZN => TL01_CLR1_n_1386);
  TL01_CLR1_g40628 : AOI211XD0BWP7T port map(A1 => TL01_CLR1_n_1194, A2 => TL01_CLR1_n_245, B => TL01_CLR1_n_1335, C => TL01_CLR1_n_1230, ZN => TL01_CLR1_n_1376);
  TL01_CLR1_g40629 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_1307, A2 => TL01_CLR1_n_690, B1 => TL01_CLR1_n_1145, B2 => TL01_CLR1_n_492, C => TL01_CLR1_n_1213, ZN => TL01_CLR1_n_1375);
  TL01_CLR1_g40630 : ND4D0BWP7T port map(A1 => TL01_CLR1_n_1316, A2 => TL01_CLR1_n_1073, A3 => TL01_CLR1_n_1207, A4 => TL01_CLR1_n_995, ZN => TL01_CLR1_n_1374);
  TL01_CLR1_g40631 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1339, A2 => TL01_CLR1_n_1304, B1 => TL01_CLR1_n_1225, B2 => vcountintern(8), ZN => TL01_CLR1_n_1373);
  TL01_CLR1_g40632 : MAOI222D1BWP7T port map(A => TL01_CLR1_n_1348, B => TL01_CLR1_n_1251, C => hcountintern(8), ZN => TL01_CLR1_n_1379);
  TL01_CLR1_g40633 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1364, A2 => TL01_CLR1_n_1119, ZN => TL01_CLR1_n_1378);
  TL01_CLR1_g40634 : MAOI222D1BWP7T port map(A => TL01_CLR1_n_1349, B => TL01_CLR1_n_1252, C => hcountintern(8), ZN => TL01_CLR1_n_1377);
  TL01_CLR1_g40635 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_1326, A2 => TL01_CLR1_n_415, B1 => TL01_CLR1_n_1098, B2 => TL01_CLR1_n_889, C1 => TL01_CLR1_n_1228, C2 => TL01_CLR1_n_430, ZN => TL01_CLR1_n_1372);
  TL01_CLR1_g40636 : OAI222D0BWP7T port map(A1 => TL01_CLR1_n_1322, A2 => TL01_CLR1_n_507, B1 => TL01_CLR1_n_315, B2 => TL01_CLR1_n_1334, C1 => TL01_CLR1_n_314, C2 => TL01_CLR1_n_1236, ZN => TL01_CLR1_n_1371);
  TL01_CLR1_g40637 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_1271, A2 => TL01_CLR1_n_735, B1 => TL01_CLR1_n_169, B2 => TL01_CLR1_n_1204, C => TL01_CLR1_n_1347, ZN => TL01_CLR1_n_1370);
  TL01_CLR1_g40638 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_1264, A2 => TL01_CLR1_n_1299, B1 => TL01_CLR1_n_1318, B2 => hcountintern(9), C1 => TL01_CLR1_n_1198, C2 => hcountintern(8), ZN => TL01_CLR1_n_1369);
  TL01_CLR1_g40639 : AOI31D0BWP7T port map(A1 => TL01_CLR1_n_1149, A2 => TL01_CLR1_n_799, A3 => TL01_CLR1_n_310, B => TL01_CLR1_n_1356, ZN => TL01_CLR1_n_1368);
  TL01_CLR1_g40640 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_880, A2 => TL01_CLR1_n_721, B1 => TL01_CLR1_n_409, B2 => TL01_CLR1_n_926, C => TL01_CLR1_n_1336, ZN => TL01_CLR1_n_1367);
  TL01_CLR1_g40641 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1337, A2 => TL01_CLR1_n_1044, B1 => TL01_CLR1_n_1031, B2 => TL01_CLR1_n_943, ZN => TL01_CLR1_n_1366);
  TL01_CLR1_g40642 : AOI211D1BWP7T port map(A1 => TL01_CLR1_n_1198, A2 => hcountintern(9), B => TL01_CLR1_n_1345, C => TL01_CLR1_n_123, ZN => TL01_CLR1_n_1365);
  TL01_CLR1_g40643 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1305, A2 => TL01_CLR1_n_1317, B1 => TL01_CLR1_n_1199, B2 => TL01_CLR1_n_166, ZN => TL01_CLR1_n_1363);
  TL01_CLR1_g40644 : AOI32D1BWP7T port map(A1 => TL01_CLR1_n_1243, A2 => TL01_CLR1_n_283, A3 => TL01_CLR1_n_313, B1 => TL01_CLR1_n_1327, B2 => TL01_CLR1_n_501, ZN => TL01_CLR1_n_1362);
  TL01_CLR1_g40645 : AOI211XD0BWP7T port map(A1 => TL01_CLR1_n_1063, A2 => TL01_CLR1_n_812, B => TL01_CLR1_n_1319, C => TL01_CLR1_n_1143, ZN => TL01_CLR1_n_1361);
  TL01_CLR1_g40646 : AOI31D0BWP7T port map(A1 => TL01_CLR1_n_1104, A2 => TL01_CLR1_n_1108, A3 => TL01_CLR1_n_562, B => TL01_CLR1_n_1338, ZN => TL01_CLR1_n_1360);
  TL01_CLR1_g40647 : AOI211XD0BWP7T port map(A1 => TL01_CLR1_n_1211, A2 => TL01_CLR1_n_1151, B => TL01_CLR1_n_1325, C => TL01_CLR1_n_1268, ZN => TL01_CLR1_n_1359);
  TL01_CLR1_g40649 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_576, A2 => TL01_CLR1_n_1303, B1 => TL01_CLR1_n_918, B2 => TL01_CLR1_n_1205, C => TL01_CLR1_n_1124, ZN => TL01_CLR1_n_1364);
  TL01_CLR1_g40650 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_1294, A2 => TL01_CLR1_n_554, B1 => TL01_CLR1_n_1158, B2 => TL01_CLR1_n_954, C1 => TL01_CLR1_n_1092, C2 => TL01_CLR1_n_928, ZN => TL01_CLR1_n_1358);
  TL01_CLR1_g40651 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_1088, A2 => TL01_CLR1_n_864, B1 => TL01_CLR1_n_1062, B2 => TL01_CLR1_n_1114, C => TL01_CLR1_n_1329, ZN => TL01_CLR1_n_1357);
  TL01_CLR1_g40652 : OAI33D1BWP7T port map(A1 => TL01_CLR1_n_379, A2 => TL01_CLR1_n_832, A3 => TL01_CLR1_n_1279, B1 => TL01_CLR1_n_368, B2 => TL01_CLR1_n_718, B3 => TL01_CLR1_n_1156, ZN => TL01_CLR1_n_1356);
  TL01_CLR1_g40653 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1321, A2 => TL01_CLR1_n_510, B1 => TL01_CLR1_n_1208, B2 => TL01_CLR1_n_579, ZN => TL01_CLR1_n_1355);
  TL01_CLR1_g40654 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1317, A2 => TL01_CLR1_n_81, B1 => TL01_CLR1_n_1199, B2 => TL01_CLR1_n_60, ZN => TL01_CLR1_n_1354);
  TL01_CLR1_g40655 : OA222D0BWP7T port map(A1 => TL01_CLR1_n_1286, A2 => TL01_CLR1_n_612, B1 => TL01_CLR1_n_931, B2 => TL01_CLR1_n_1088, C1 => TL01_CLR1_n_919, C2 => TL01_CLR1_n_1153, Z => TL01_CLR1_n_1353);
  TL01_CLR1_g40656 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_1180, A2 => TL01_CLR1_n_1157, B1 => TL01_CLR1_n_1300, B2 => TL01_CLR1_n_831, C1 => TL01_CLR1_n_1149, C2 => TL01_CLR1_n_786, ZN => TL01_CLR1_n_1352);
  TL01_CLR1_g40657 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1315, A2 => TL01_CLR1_n_283, ZN => TL01_CLR1_n_1350);
  TL01_CLR1_g40658 : OAI31D0BWP7T port map(A1 => TL01_CLR1_n_599, A2 => TL01_CLR1_n_867, A3 => TL01_CLR1_n_1249, B => TL01_CLR1_n_1312, ZN => TL01_CLR1_n_1349);
  TL01_CLR1_g40659 : OAI31D0BWP7T port map(A1 => TL01_CLR1_n_585, A2 => TL01_CLR1_n_866, A3 => TL01_CLR1_n_1248, B => TL01_CLR1_n_1311, ZN => TL01_CLR1_n_1348);
  TL01_CLR1_g40660 : OA33D0BWP7T port map(A1 => vcountintern(4), A2 => TL01_CLR1_n_386, A3 => TL01_CLR1_n_1271, B1 => vcountintern(5), B2 => TL01_CLR1_n_1019, B3 => TL01_CLR1_n_1165, Z => TL01_CLR1_n_1347);
  TL01_CLR1_g40661 : OAI31D0BWP7T port map(A1 => vcountintern(4), A2 => TL01_CLR1_n_384, A3 => TL01_CLR1_n_1272, B => TL01_CLR1_n_1262, ZN => TL01_CLR1_n_1346);
  TL01_CLR1_g40662 : OA21D0BWP7T port map(A1 => TL01_CLR1_n_1198, A2 => TL01_CLR1_n_165, B => TL01_CLR1_n_1318, Z => TL01_CLR1_n_1345);
  TL01_CLR1_g40663 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_1005, A2 => TL01_CLR1_n_1150, B => TL01_CLR1_n_1278, C => TL01_CLR1_n_1285, ZN => TL01_CLR1_n_1344);
  TL01_CLR1_g40664 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_1151, A2 => TL01_CLR1_n_949, B1 => TL01_CLR1_n_1218, B2 => TL01_CLR1_n_821, C => TL01_CLR1_n_1328, ZN => TL01_CLR1_n_1343);
  TL01_CLR1_g40665 : AOI31D0BWP7T port map(A1 => TL01_CLR1_n_1233, A2 => TL01_CLR1_n_430, A3 => TL01_CLR1_n_283, B => TL01_CLR1_n_1240, ZN => TL01_CLR1_n_1342);
  TL01_CLR1_g40666 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_744, A2 => TL01_CLR1_n_571, B1 => TL01_CLR1_n_498, B2 => TL01_CLR1_n_922, C => TL01_CLR1_n_1314, ZN => TL01_CLR1_n_1351);
  TL01_CLR1_g40667 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1273, A2 => TL01_CLR1_n_48, B1 => TL01_CLR1_n_1244, B2 => TL01_CLR1_n_742, ZN => TL01_CLR1_n_1340);
  TL01_CLR1_g40668 : OAI32D1BWP7T port map(A1 => TL01_CLR1_n_176, A2 => TL01_CLR1_n_891, A3 => TL01_CLR1_n_1250, B1 => TL01_CLR1_n_107, B2 => TL01_CLR1_n_1253, ZN => TL01_CLR1_n_1339);
  TL01_CLR1_g40669 : OAI32D1BWP7T port map(A1 => TL01_CLR1_n_312, A2 => TL01_CLR1_n_387, A3 => TL01_CLR1_n_1242, B1 => TL01_CLR1_n_847, B2 => TL01_CLR1_n_1101, ZN => TL01_CLR1_n_1338);
  TL01_CLR1_g40670 : OAI222D0BWP7T port map(A1 => TL01_CLR1_n_1269, A2 => TL01_CLR1_n_375, B1 => TL01_CLR1_n_745, B2 => TL01_CLR1_n_1195, C1 => TL01_CLR1_n_694, C2 => TL01_CLR1_n_718, ZN => TL01_CLR1_n_1337);
  TL01_CLR1_g40671 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_1260, A2 => TL01_CLR1_n_410, B1 => TL01_CLR1_n_1074, B2 => TL01_CLR1_n_751, C1 => TL01_CLR1_n_817, C2 => TL01_CLR1_n_816, ZN => TL01_CLR1_n_1336);
  TL01_CLR1_g40672 : OAI31D0BWP7T port map(A1 => TL01_CLR1_n_373, A2 => TL01_CLR1_n_1105, A3 => TL01_CLR1_n_1220, B => TL01_CLR1_n_1324, ZN => TL01_CLR1_n_1335);
  TL01_CLR1_g40673 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1287, A2 => TL01_CLR1_n_719, B1 => TL01_CLR1_n_1280, B2 => TL01_CLR1_n_831, ZN => TL01_CLR1_n_1334);
  TL01_CLR1_g40674 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_1224, A2 => FE_PHN123_char2posx_8, B1 => TL01_CLR1_n_1224, B2 => FE_PHN123_char2posx_8, ZN => TL01_CLR1_n_1333);
  TL01_CLR1_g40675 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_1306, A2 => TL01_CLR1_n_805, B1 => TL01_CLR1_n_1223, B2 => TL01_CLR1_n_976, ZN => TL01_CLR1_n_1332);
  TL01_CLR1_g40676 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_1221, A2 => char1posx(8), B1 => TL01_CLR1_n_1221, B2 => char1posx(8), ZN => TL01_CLR1_n_1331);
  TL01_CLR1_g40677 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_662, A2 => TL01_CLR1_n_1061, B1 => TL01_CLR1_n_1011, B2 => TL01_CLR1_n_1289, ZN => TL01_CLR1_n_1341);
  TL01_CLR1_g40678 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_712, A2 => TL01_CLR1_n_1099, B => TL01_CLR1_n_1239, C => TL01_CLR1_n_1215, ZN => TL01_CLR1_n_1330);
  TL01_CLR1_g40679 : OA31D1BWP7T port map(A1 => TL01_CLR1_n_237, A2 => TL01_CLR1_n_1106, A3 => TL01_CLR1_n_1220, B => TL01_CLR1_n_1130, Z => TL01_CLR1_n_1329);
  TL01_CLR1_g40680 : IAO21D0BWP7T port map(A1 => TL01_CLR1_n_684, A2 => TL01_CLR1_n_310, B => TL01_CLR1_n_1288, ZN => TL01_CLR1_n_1328);
  TL01_CLR1_g40681 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_1197, A2 => TL01_CLR1_n_1107, B1 => TL01_CLR1_n_1029, B2 => TL01_CLR1_n_1094, C => TL01_CLR1_n_1181, ZN => TL01_CLR1_n_1327);
  TL01_CLR1_g40682 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_1080, A2 => TL01_CLR1_n_1077, B1 => TL01_CLR1_n_962, B2 => TL01_CLR1_n_972, C => TL01_CLR1_n_1275, ZN => TL01_CLR1_n_1326);
  TL01_CLR1_g40683 : OAI31D0BWP7T port map(A1 => TL01_CLR1_n_309, A2 => TL01_CLR1_n_1161, A3 => TL01_CLR1_n_1220, B => TL01_CLR1_n_1231, ZN => TL01_CLR1_n_1325);
  TL01_CLR1_g40684 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1261, A2 => TL01_CLR1_n_1098, B1 => TL01_CLR1_n_1116, B2 => TL01_CLR1_n_1022, ZN => TL01_CLR1_n_1324);
  TL01_CLR1_g40685 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1123, A2 => TL01_CLR1_n_1188, B1 => TL01_CLR1_n_1254, B2 => TL01_CLR1_n_158, ZN => TL01_CLR1_n_1323);
  TL01_CLR1_g40686 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_1196, A2 => TL01_CLR1_n_1160, B1 => TL01_CLR1_n_1162, B2 => TL01_CLR1_n_1076, C => TL01_CLR1_n_1234, ZN => TL01_CLR1_n_1322);
  TL01_CLR1_g40687 : AO221D0BWP7T port map(A1 => TL01_CLR1_n_1042, A2 => TL01_CLR1_n_1076, B1 => TL01_CLR1_n_977, B2 => TL01_CLR1_n_961, C => TL01_CLR1_n_1274, Z => TL01_CLR1_n_1321);
  TL01_CLR1_g40688 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_1247, A2 => TL01_CLR1_n_840, B => TL01_CLR1_n_1116, ZN => TL01_CLR1_n_1320);
  TL01_CLR1_g40689 : OAI32D1BWP7T port map(A1 => TL01_CLR1_n_723, A2 => TL01_CLR1_n_1040, A3 => TL01_CLR1_n_1220, B1 => TL01_CLR1_n_1036, B2 => TL01_CLR1_n_1217, ZN => TL01_CLR1_n_1319);
  TL01_CLR1_g40690 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_1247, A2 => TL01_CLR1_n_42, B1 => TL01_CLR1_n_957, B2 => TL01_CLR1_n_751, C1 => TL01_CLR1_n_817, C2 => TL01_CLR1_n_736, ZN => TL01_CLR1_n_1316);
  TL01_CLR1_g40691 : OAI31D0BWP7T port map(A1 => TL01_CLR1_n_103, A2 => TL01_CLR1_n_558, A3 => TL01_CLR1_n_1103, B => TL01_CLR1_n_1302, ZN => TL01_CLR1_n_1315);
  TL01_CLR1_g40692 : AOI211XD0BWP7T port map(A1 => TL01_CLR1_n_677, A2 => TL01_CLR1_n_574, B => TL01_CLR1_n_1267, C => TL01_CLR1_n_790, ZN => TL01_CLR1_n_1314);
  TL01_CLR1_g40693 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_1238, A2 => TL01_CLR1_n_642, B1 => TL01_CLR1_n_1031, B2 => TL01_CLR1_n_857, C1 => TL01_CLR1_n_1095, C2 => TL01_CLR1_n_742, ZN => TL01_CLR1_n_1313);
  TL01_CLR1_g40694 : OA221D0BWP7T port map(A1 => TL01_CLR1_n_1249, A2 => TL01_CLR1_n_862, B1 => TL01_CLR1_n_158, B2 => TL01_CLR1_n_1045, C => TL01_CLR1_n_1182, Z => TL01_CLR1_n_1312);
  TL01_CLR1_g40695 : OA221D0BWP7T port map(A1 => TL01_CLR1_n_1248, A2 => TL01_CLR1_n_861, B1 => TL01_CLR1_n_158, B2 => TL01_CLR1_n_1053, C => TL01_CLR1_n_1193, Z => TL01_CLR1_n_1311);
  TL01_CLR1_g40696 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_755, A2 => TL01_CLR1_n_946, B => TL01_CLR1_n_1259, C => TL01_CLR1_n_1007, ZN => TL01_CLR1_n_1310);
  TL01_CLR1_g40697 : AOI33D1BWP7T port map(A1 => TL01_CLR1_n_1189, A2 => TL01_CLR1_n_579, A3 => TL01_CLR1_n_311, B1 => TL01_CLR1_n_1104, B2 => TL01_CLR1_n_1042, B3 => TL01_CLR1_n_565, ZN => TL01_CLR1_n_1309);
  TL01_CLR1_g40698 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_717, A2 => TL01_CLR1_n_324, B1 => TL01_CLR1_n_1269, B2 => TL01_CLR1_n_385, ZN => TL01_CLR1_n_1308);
  TL01_CLR1_g40699 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1269, A2 => TL01_CLR1_n_388, B1 => TL01_CLR1_n_718, B2 => TL01_CLR1_n_247, ZN => TL01_CLR1_n_1307);
  TL01_CLR1_g40700 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_1169, A2 => char1posx(8), B1 => TL01_CLR1_n_1169, B2 => char1posx(8), ZN => TL01_CLR1_n_1318);
  TL01_CLR1_g40701 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_1166, A2 => FE_PHN123_char2posx_8, B1 => TL01_CLR1_n_1166, B2 => FE_PHN123_char2posx_8, ZN => TL01_CLR1_n_1317);
  TL01_CLR1_g40702 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_1199, A2 => TL01_CLR1_n_81, Z => TL01_CLR1_n_1305);
  TL01_CLR1_g40703 : NR3D0BWP7T port map(A1 => TL01_CLR1_n_1250, A2 => TL01_CLR1_n_664, A3 => TL01_CLR1_n_871, ZN => TL01_CLR1_n_1304);
  TL01_CLR1_g40704 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_1070, A2 => TL01_CLR1_n_849, B1 => TL01_CLR1_n_1109, B2 => TL01_CLR1_n_72, C => TL01_CLR1_n_1258, ZN => TL01_CLR1_n_1303);
  TL01_CLR1_g40705 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_1178, A2 => TL01_CLR1_n_1177, B => TL01_CLR1_n_245, ZN => TL01_CLR1_n_1302);
  TL01_CLR1_g40706 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_1171, A2 => vcountintern(7), B1 => vcountintern(6), B2 => TL01_CLR1_n_914, C => TL01_CLR1_n_1008, ZN => TL01_CLR1_n_1301);
  TL01_CLR1_g40707 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_1161, A2 => TL01_CLR1_n_820, B1 => TL01_CLR1_n_680, B2 => TL01_CLR1_n_1038, C => TL01_CLR1_n_1229, ZN => TL01_CLR1_n_1300);
  TL01_CLR1_g40708 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_153, A2 => TL01_CLR1_n_1014, B => TL01_CLR1_n_1201, C => TL01_CLR1_n_158, ZN => TL01_CLR1_n_1299);
  TL01_CLR1_g40709 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_1171, A2 => TL01_CLR1_n_1020, B1 => vcountintern(7), B2 => TL01_CLR1_n_914, C => TL01_CLR1_n_106, ZN => TL01_CLR1_n_1298);
  TL01_CLR1_g40710 : OA21D0BWP7T port map(A1 => TL01_CLR1_n_1153, A2 => TL01_CLR1_n_686, B => TL01_CLR1_n_1266, Z => TL01_CLR1_n_1297);
  TL01_CLR1_g40711 : AOI32D1BWP7T port map(A1 => TL01_CLR1_n_1104, A2 => TL01_CLR1_n_1162, A3 => TL01_CLR1_n_684, B1 => TL01_CLR1_n_1024, B2 => TL01_CLR1_n_1149, ZN => TL01_CLR1_n_1296);
  TL01_CLR1_g40712 : AOI211D0BWP7T port map(A1 => TL01_CLR1_n_384, A2 => vcountintern(4), B => TL01_CLR1_n_1272, C => TL01_CLR1_n_701, ZN => TL01_CLR1_n_1295);
  TL01_CLR1_g40713 : OAI31D0BWP7T port map(A1 => char1perc(0), A2 => TL01_CLR1_n_623, A3 => TL01_CLR1_n_1039, B => TL01_CLR1_n_1235, ZN => TL01_CLR1_n_1294);
  TL01_CLR1_g40714 : IOA21D0BWP7T port map(A1 => TL01_CLR1_n_1227, A2 => TL01_CLR1_n_68, B => TL01_CLR1_n_147, ZN => TL01_CLR1_n_1293);
  TL01_CLR1_g40715 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1210, A2 => vcountintern(8), B1 => TL01_CLR1_n_1163, B2 => vcountintern(9), ZN => TL01_CLR1_n_1292);
  TL01_CLR1_g40716 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_1225, A2 => vcountintern(9), B => TL01_CLR1_n_147, ZN => TL01_CLR1_n_1291);
  TL01_CLR1_g40717 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_1185, A2 => TL01_CLR1_n_489, A3 => TL01_CLR1_n_311, ZN => TL01_CLR1_n_1290);
  TL01_CLR1_g40718 : NR4D0BWP7T port map(A1 => TL01_CLR1_n_1132, A2 => TL01_CLR1_n_1168, A3 => TL01_CLR1_n_930, A4 => TL01_CLR1_n_843, ZN => TL01_CLR1_n_1306);
  TL01_CLR1_g40719 : AOI32D1BWP7T port map(A1 => TL01_CLR1_n_728, A2 => TL01_CLR1_n_566, A3 => TL01_CLR1_n_71, B1 => TL01_CLR1_n_827, B2 => TL01_CLR1_n_1191, ZN => TL01_CLR1_n_1289);
  TL01_CLR1_g40720 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_1136, A2 => TL01_CLR1_n_727, B1 => TL01_CLR1_n_1151, B2 => TL01_CLR1_n_622, C1 => TL01_CLR1_n_1157, C2 => TL01_CLR1_n_1028, ZN => TL01_CLR1_n_1288);
  TL01_CLR1_g40721 : OAI222D0BWP7T port map(A1 => TL01_CLR1_n_1159, A2 => TL01_CLR1_n_822, B1 => TL01_CLR1_n_739, B2 => TL01_CLR1_n_1155, C1 => TL01_CLR1_n_674, C2 => TL01_CLR1_n_1038, ZN => TL01_CLR1_n_1287);
  TL01_CLR1_g40722 : OA21D0BWP7T port map(A1 => TL01_CLR1_n_1101, A2 => TL01_CLR1_n_1029, B => TL01_CLR1_n_1232, Z => TL01_CLR1_n_1286);
  TL01_CLR1_g40723 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_1218, A2 => TL01_CLR1_n_819, B1 => TL01_CLR1_n_1151, B2 => TL01_CLR1_n_850, C1 => TL01_CLR1_n_1149, C2 => TL01_CLR1_n_870, ZN => TL01_CLR1_n_1285);
  TL01_CLR1_g40724 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1175, A2 => TL01_CLR1_n_313, B1 => TL01_CLR1_n_1139, B2 => TL01_CLR1_n_1099, ZN => TL01_CLR1_n_1284);
  TL01_CLR1_g40725 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_1158, A2 => TL01_CLR1_n_898, B1 => TL01_CLR1_n_1092, B2 => TL01_CLR1_n_651, C1 => TL01_CLR1_n_1092, C2 => TL01_CLR1_n_1026, ZN => TL01_CLR1_n_1283);
  TL01_CLR1_g40726 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_811, A2 => TL01_CLR1_n_713, B1 => TL01_CLR1_n_755, B2 => TL01_CLR1_n_1072, C => TL01_CLR1_n_1186, ZN => TL01_CLR1_n_1282);
  TL01_CLR1_g40727 : OA22D0BWP7T port map(A1 => TL01_CLR1_n_1146, A2 => TL01_CLR1_n_1088, B1 => TL01_CLR1_n_1101, B2 => TL01_CLR1_n_1173, Z => TL01_CLR1_n_1281);
  TL01_CLR1_g40728 : OAI222D0BWP7T port map(A1 => TL01_CLR1_n_1156, A2 => TL01_CLR1_n_680, B1 => TL01_CLR1_n_726, B2 => TL01_CLR1_n_910, C1 => TL01_CLR1_n_558, C2 => TL01_CLR1_n_1155, ZN => TL01_CLR1_n_1280);
  TL01_CLR1_g40729 : AOI32D1BWP7T port map(A1 => TL01_CLR1_n_1157, A2 => TL01_CLR1_n_740, A3 => TL01_CLR1_n_233, B1 => TL01_CLR1_n_1160, B2 => TL01_CLR1_n_557, ZN => TL01_CLR1_n_1279);
  TL01_CLR1_g40730 : AOI32D1BWP7T port map(A1 => TL01_CLR1_n_1162, A2 => TL01_CLR1_n_719, A3 => TL01_CLR1_n_620, B1 => TL01_CLR1_n_1218, B2 => TL01_CLR1_n_902, ZN => TL01_CLR1_n_1278);
  TL01_CLR1_g40731 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_378, A2 => TL01_CLR1_n_1059, B1 => TL01_CLR1_n_378, B2 => TL01_CLR1_n_1216, ZN => TL01_CLR1_n_1277);
  TL01_CLR1_g40732 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_1214, A2 => TL01_CLR1_n_1149, B1 => TL01_CLR1_n_1219, B2 => TL01_CLR1_n_908, ZN => TL01_CLR1_n_1276);
  TL01_CLR1_g40733 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_45, A2 => TL01_CLR1_n_1028, B1 => TL01_CLR1_n_1197, B2 => TL01_CLR1_n_1103, ZN => TL01_CLR1_n_1275);
  TL01_CLR1_g40734 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1197, A2 => TL01_CLR1_n_1041, B1 => TL01_CLR1_n_1029, B2 => TL01_CLR1_n_1035, ZN => TL01_CLR1_n_1274);
  TL01_CLR1_g40735 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1195, A2 => TL01_CLR1_n_513, B1 => TL01_CLR1_n_718, B2 => TL01_CLR1_n_572, ZN => TL01_CLR1_n_1273);
  TL01_CLR1_g40736 : NR3D0BWP7T port map(A1 => TL01_CLR1_n_1161, A2 => TL01_CLR1_n_883, A3 => TL01_CLR1_n_683, ZN => TL01_CLR1_n_1268);
  TL01_CLR1_g40737 : OAI211D1BWP7T port map(A1 => vcountintern(0), A2 => TL01_CLR1_n_797, B => TL01_CLR1_n_1023, C => TL01_CLR1_n_1134, ZN => TL01_CLR1_n_1267);
  TL01_CLR1_g40738 : OAI31D0BWP7T port map(A1 => TL01_CLR1_n_825, A2 => TL01_CLR1_n_1057, A3 => TL01_CLR1_n_1115, B => TL01_CLR1_n_1100, ZN => TL01_CLR1_n_1266);
  TL01_CLR1_g40739 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_929, A2 => TL01_CLR1_n_750, B1 => TL01_CLR1_n_747, B2 => TL01_CLR1_n_818, C => TL01_CLR1_n_1209, ZN => TL01_CLR1_n_1265);
  TL01_CLR1_g40740 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1190, A2 => TL01_CLR1_n_1187, ZN => TL01_CLR1_n_1264);
  TL01_CLR1_g40741 : OA221D0BWP7T port map(A1 => TL01_CLR1_n_1106, A2 => TL01_CLR1_n_820, B1 => TL01_CLR1_n_600, B2 => TL01_CLR1_n_1094, C => TL01_CLR1_n_1184, Z => TL01_CLR1_n_1263);
  TL01_CLR1_g40742 : ND4D0BWP7T port map(A1 => TL01_CLR1_n_1164, A2 => TL01_CLR1_n_982, A3 => TL01_CLR1_n_606, A4 => TL01_CLR1_n_86, ZN => TL01_CLR1_n_1262);
  TL01_CLR1_g40743 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_1122, A2 => TL01_CLR1_n_951, A3 => TL01_CLR1_n_836, ZN => TL01_CLR1_n_1261);
  TL01_CLR1_g40744 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_508, A2 => TL01_CLR1_n_600, B => TL01_CLR1_n_1144, C => TL01_CLR1_n_951, ZN => TL01_CLR1_n_1260);
  TL01_CLR1_g40745 : OAI31D0BWP7T port map(A1 => TL01_CLR1_n_698, A2 => TL01_CLR1_n_1069, A3 => TL01_CLR1_n_1115, B => TL01_CLR1_n_492, ZN => TL01_CLR1_n_1259);
  TL01_CLR1_g40746 : OAI31D0BWP7T port map(A1 => TL01_CLR1_n_456, A2 => TL01_CLR1_n_661, A3 => TL01_CLR1_n_1009, B => TL01_CLR1_n_1203, ZN => TL01_CLR1_n_1258);
  TL01_CLR1_g40747 : AOI31D0BWP7T port map(A1 => TL01_CLR1_n_455, A2 => TL01_CLR1_char1_sprite_sprite_0, A3 => TL01_CLR1_n_1084, B => TL01_CLR1_n_1192, ZN => TL01_CLR1_n_1257);
  TL01_CLR1_g40748 : AOI211D0BWP7T port map(A1 => TL01_CLR1_n_803, A2 => vcountintern(7), B => TL01_CLR1_n_1126, C => TL01_CLR1_n_169, ZN => TL01_CLR1_n_1256);
  TL01_CLR1_g40749 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1142, A2 => TL01_CLR1_n_1031, B1 => TL01_CLR1_n_1095, B2 => TL01_CLR1_n_953, ZN => TL01_CLR1_n_1255);
  TL01_CLR1_g40750 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1141, A2 => TL01_CLR1_n_807, B1 => TL01_CLR1_n_1012, B2 => hcountintern(7), ZN => TL01_CLR1_n_1254);
  TL01_CLR1_g40751 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1027, A2 => TL01_CLR1_n_1172, B1 => TL01_CLR1_n_913, B2 => TL01_CLR1_n_169, ZN => TL01_CLR1_n_1253);
  TL01_CLR1_g40752 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_86, A2 => TL01_CLR1_n_606, B => TL01_CLR1_n_1164, C => TL01_CLR1_n_982, ZN => TL01_CLR1_n_1272);
  TL01_CLR1_g40753 : AO211D0BWP7T port map(A1 => TL01_CLR1_n_603, A2 => vcountintern(5), B => TL01_CLR1_n_1165, C => TL01_CLR1_n_980, Z => TL01_CLR1_n_1271);
  TL01_CLR1_g40754 : INR2D1BWP7T port map(A1 => TL01_CLR1_n_1223, B1 => TL01_CLR1_n_976, ZN => TL01_CLR1_n_1270);
  TL01_CLR1_g40755 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_1055, A2 => char2posx(7), B => TL01_CLR1_n_1224, ZN => TL01_CLR1_n_1252);
  TL01_CLR1_g40756 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_1054, A2 => char1posx(7), B => TL01_CLR1_n_1221, ZN => TL01_CLR1_n_1251);
  TL01_CLR1_g40757 : CKAN2D1BWP7T port map(A1 => TL01_CLR1_n_1195, A2 => TL01_CLR1_n_718, Z => TL01_CLR1_n_1269);
  TL01_CLR1_g40758 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1088, A2 => TL01_CLR1_n_1001, B1 => TL01_CLR1_n_1153, B2 => TL01_CLR1_n_903, ZN => TL01_CLR1_n_1245);
  TL01_CLR1_g40759 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_1150, A2 => TL01_CLR1_n_233, B => TL01_CLR1_n_1219, ZN => TL01_CLR1_n_1244);
  TL01_CLR1_g40760 : OAI222D0BWP7T port map(A1 => TL01_CLR1_n_1094, A2 => TL01_CLR1_n_739, B1 => TL01_CLR1_n_822, B2 => TL01_CLR1_n_1107, C1 => TL01_CLR1_n_674, C2 => TL01_CLR1_n_830, ZN => TL01_CLR1_n_1243);
  TL01_CLR1_g40761 : OA222D0BWP7T port map(A1 => TL01_CLR1_n_1101, A2 => TL01_CLR1_n_877, B1 => TL01_CLR1_n_558, B2 => TL01_CLR1_n_1094, C1 => TL01_CLR1_n_730, C2 => TL01_CLR1_n_910, Z => TL01_CLR1_n_1242);
  TL01_CLR1_g40762 : AOI32D1BWP7T port map(A1 => TL01_CLR1_n_1089, A2 => TL01_CLR1_n_45, A3 => TL01_CLR1_n_307, B1 => TL01_CLR1_n_1098, B2 => TL01_CLR1_n_998, ZN => TL01_CLR1_n_1241);
  TL01_CLR1_g40763 : AO21D0BWP7T port map(A1 => TL01_CLR1_n_1102, A2 => TL01_CLR1_n_939, B => TL01_CLR1_n_1206, Z => TL01_CLR1_n_1240);
  TL01_CLR1_g40764 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1152, A2 => TL01_CLR1_n_819, B1 => TL01_CLR1_n_1087, B2 => TL01_CLR1_n_851, ZN => TL01_CLR1_n_1239);
  TL01_CLR1_g40765 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1127, A2 => TL01_CLR1_n_601, B1 => TL01_CLR1_n_1029, B2 => TL01_CLR1_n_1037, ZN => TL01_CLR1_n_1238);
  TL01_CLR1_g40766 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1158, A2 => TL01_CLR1_n_819, B1 => TL01_CLR1_n_1138, B2 => TL01_CLR1_n_682, ZN => TL01_CLR1_n_1237);
  TL01_CLR1_g40767 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1089, A2 => TL01_CLR1_n_1154, B1 => TL01_CLR1_n_1149, B2 => TL01_CLR1_n_675, ZN => TL01_CLR1_n_1236);
  TL01_CLR1_g40768 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1102, A2 => TL01_CLR1_n_1028, B1 => TL01_CLR1_n_1133, B2 => TL01_CLR1_n_904, ZN => TL01_CLR1_n_1235);
  TL01_CLR1_g40769 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1155, A2 => TL01_CLR1_n_1029, B1 => TL01_CLR1_n_962, B2 => TL01_CLR1_n_1038, ZN => TL01_CLR1_n_1234);
  TL01_CLR1_g40770 : AO21D0BWP7T port map(A1 => TL01_CLR1_n_45, A2 => TL01_CLR1_n_557, B => TL01_CLR1_n_1183, Z => TL01_CLR1_n_1233);
  TL01_CLR1_g40771 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_1135, A2 => TL01_CLR1_n_731, B1 => TL01_CLR1_n_1088, B2 => TL01_CLR1_n_623, ZN => TL01_CLR1_n_1232);
  TL01_CLR1_g40772 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_48, A2 => TL01_CLR1_n_948, B1 => TL01_CLR1_n_1149, B2 => TL01_CLR1_n_865, ZN => TL01_CLR1_n_1231);
  TL01_CLR1_g40773 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_1091, A2 => TL01_CLR1_n_991, B1 => TL01_CLR1_n_1158, B2 => TL01_CLR1_n_902, ZN => TL01_CLR1_n_1230);
  TL01_CLR1_g40774 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_1160, A2 => TL01_CLR1_n_814, B1 => TL01_CLR1_n_1155, B2 => TL01_CLR1_n_600, ZN => TL01_CLR1_n_1229);
  TL01_CLR1_g40775 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_1131, A2 => TL01_CLR1_n_822, B1 => TL01_CLR1_n_45, B2 => TL01_CLR1_n_740, ZN => TL01_CLR1_n_1228);
  TL01_CLR1_g40776 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1172, A2 => vcountintern(7), B1 => TL01_CLR1_n_913, B2 => vcountintern(6), ZN => TL01_CLR1_n_1250);
  TL01_CLR1_g40777 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1083, A2 => hcountintern(7), B1 => TL01_CLR1_n_917, B2 => hcountintern(6), ZN => TL01_CLR1_n_1249);
  TL01_CLR1_g40778 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1082, A2 => hcountintern(7), B1 => TL01_CLR1_n_920, B2 => hcountintern(6), ZN => TL01_CLR1_n_1248);
  TL01_CLR1_g40779 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_368, A2 => TL01_CLR1_n_319, B => TL01_CLR1_n_1195, ZN => TL01_CLR1_n_1247);
  TL01_CLR1_g40780 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1140, A2 => TL01_CLR1_n_1013, B1 => TL01_CLR1_n_915, B2 => TL01_CLR1_n_769, ZN => TL01_CLR1_n_1246);
  TL01_CLR1_g40781 : INVD1BWP7T port map(I => TL01_CLR1_n_1219, ZN => TL01_CLR1_n_1218);
  TL01_CLR1_g40782 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_1033, A2 => TL01_CLR1_n_316, B1 => TL01_CLR1_n_620, B2 => TL01_CLR1_n_722, C => TL01_CLR1_n_947, ZN => TL01_CLR1_n_1217);
  TL01_CLR1_g40783 : OAI32D1BWP7T port map(A1 => TL01_CLR1_n_934, A2 => TL01_CLR1_n_848, A3 => TL01_CLR1_n_1011, B1 => orientationp2, B2 => TL01_CLR1_n_1086, ZN => TL01_CLR1_n_1216);
  TL01_CLR1_g40784 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_1108, A2 => TL01_CLR1_n_620, A3 => TL01_CLR1_n_283, ZN => TL01_CLR1_n_1215);
  TL01_CLR1_g40785 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_723, A2 => TL01_CLR1_n_1032, B => TL01_CLR1_n_1066, C => TL01_CLR1_n_782, ZN => TL01_CLR1_n_1214);
  TL01_CLR1_g40786 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_755, A2 => TL01_CLR1_n_860, B => TL01_CLR1_n_897, C => TL01_CLR1_n_1129, ZN => TL01_CLR1_n_1213);
  TL01_CLR1_g40787 : ND4D0BWP7T port map(A1 => TL01_CLR1_n_1044, A2 => TL01_CLR1_n_752, A3 => TL01_CLR1_n_582, A4 => TL01_CLR1_n_238, ZN => TL01_CLR1_n_1212);
  TL01_CLR1_g40788 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_306, A2 => TL01_CLR1_n_724, B => TL01_CLR1_n_1058, C => TL01_CLR1_n_773, ZN => TL01_CLR1_n_1211);
  TL01_CLR1_g40789 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_1170, B1 => TL01_CLR1_n_1163, ZN => TL01_CLR1_n_1210);
  TL01_CLR1_g40790 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_956, A2 => TL01_CLR1_n_751, B1 => TL01_CLR1_n_952, B2 => TL01_CLR1_n_682, C => TL01_CLR1_n_1121, ZN => TL01_CLR1_n_1209);
  TL01_CLR1_g40791 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_1040, A2 => TL01_CLR1_n_820, B1 => TL01_CLR1_n_600, B2 => TL01_CLR1_n_1035, C => TL01_CLR1_n_1117, ZN => TL01_CLR1_n_1208);
  TL01_CLR1_g40792 : IND3D1BWP7T port map(A1 => TL01_CLR1_n_508, B1 => TL01_CLR1_n_402, B2 => TL01_CLR1_n_1056, ZN => TL01_CLR1_n_1207);
  TL01_CLR1_g40793 : INR3D0BWP7T port map(A1 => TL01_CLR1_n_1104, B1 => TL01_CLR1_n_493, B2 => TL01_CLR1_n_1080, ZN => TL01_CLR1_n_1206);
  TL01_CLR1_g40794 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_1060, A2 => orientationp1, B => TL01_CLR1_n_1071, ZN => TL01_CLR1_n_1205);
  TL01_CLR1_g40795 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_958, A2 => TL01_CLR1_n_1016, B1 => TL01_CLR1_n_804, B2 => TL01_CLR1_n_107, ZN => TL01_CLR1_n_1204);
  TL01_CLR1_g40796 : IOA21D0BWP7T port map(A1 => TL01_CLR1_n_1109, A2 => TL01_CLR1_n_455, B => orientationp1, ZN => TL01_CLR1_n_1203);
  TL01_CLR1_g40797 : AOI211D1BWP7T port map(A1 => TL01_CLR1_n_502, A2 => TL01_CLR1_n_326, B => TL01_CLR1_n_1106, C => TL01_CLR1_n_683, ZN => TL01_CLR1_n_1202);
  TL01_CLR1_g40798 : IOA21D1BWP7T port map(A1 => TL01_CLR1_n_1014, A2 => TL01_CLR1_n_82, B => TL01_CLR1_n_809, ZN => TL01_CLR1_n_1201);
  TL01_CLR1_g40799 : INR2XD0BWP7T port map(A1 => char2posy(7), B1 => TL01_CLR1_n_1147, ZN => TL01_CLR1_n_1227);
  TL01_CLR1_g40800 : AOI211XD0BWP7T port map(A1 => TL01_CLR1_n_1011, A2 => TL01_CLR1_n_566, B => TL01_CLR1_n_827, C => TL01_CLR1_n_986, ZN => TL01_CLR1_n_1226);
  TL01_CLR1_g40801 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_1148, B1 => char1posy(7), ZN => TL01_CLR1_n_1225);
  TL01_CLR1_g40802 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1055, A2 => char2posx(7), ZN => TL01_CLR1_n_1224);
  TL01_CLR1_g40803 : IND3D1BWP7T port map(A1 => TL01_CLR1_n_1168, B1 => TL01_CLR1_n_944, B2 => TL01_CLR1_n_997, ZN => TL01_CLR1_n_1223);
  TL01_CLR1_g40804 : INR2XD0BWP7T port map(A1 => TL01_CLR1_n_1013, B1 => TL01_CLR1_n_1140, ZN => TL01_CLR1_n_1222);
  TL01_CLR1_g40805 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1054, A2 => char1posx(7), ZN => TL01_CLR1_n_1221);
  TL01_CLR1_g40806 : NR3D0BWP7T port map(A1 => TL01_CLR1_n_1081, A2 => TL01_CLR1_n_812, A3 => TL01_CLR1_n_752, ZN => TL01_CLR1_n_1220);
  TL01_CLR1_g40807 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1151, A2 => TL01_CLR1_n_684, ZN => TL01_CLR1_n_1219);
  TL01_CLR1_g40808 : INVD0BWP7T port map(I => TL01_CLR1_n_1197, ZN => TL01_CLR1_n_1196);
  TL01_CLR1_g40809 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1097, A2 => TL01_CLR1_n_600, B1 => TL01_CLR1_n_1080, B2 => TL01_CLR1_n_621, ZN => TL01_CLR1_n_1194);
  TL01_CLR1_g40810 : IOA21D1BWP7T port map(A1 => TL01_CLR1_n_1053, A2 => TL01_CLR1_n_82, B => TL01_CLR1_n_1082, ZN => TL01_CLR1_n_1193);
  TL01_CLR1_g40811 : OAI32D1BWP7T port map(A1 => TL01_CLR1_n_911, A2 => TL01_CLR1_char1_sprite_sprite_0, A3 => TL01_CLR1_n_1009, B1 => TL01_CLR1_n_1085, B2 => TL01_CLR1_n_661, ZN => TL01_CLR1_n_1192);
  TL01_CLR1_g40812 : OAI32D1BWP7T port map(A1 => TL01_CLR1_n_924, A2 => TL01_CLR1_n_1003, A3 => TL01_CLR1_n_516, B1 => TL01_CLR1_n_970, B2 => TL01_CLR1_n_378, ZN => TL01_CLR1_n_1191);
  TL01_CLR1_g40813 : MAOI222D1BWP7T port map(A => TL01_CLR1_n_984, B => TL01_CLR1_n_616, C => hcountintern(5), ZN => TL01_CLR1_n_1190);
  TL01_CLR1_g40814 : OAI222D0BWP7T port map(A1 => TL01_CLR1_n_1037, A2 => TL01_CLR1_n_680, B1 => TL01_CLR1_n_601, B2 => TL01_CLR1_n_910, C1 => TL01_CLR1_n_558, C2 => TL01_CLR1_n_1035, ZN => TL01_CLR1_n_1189);
  TL01_CLR1_g40815 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1012, A2 => hcountintern(7), B1 => TL01_CLR1_n_807, B2 => hcountintern(6), ZN => TL01_CLR1_n_1188);
  TL01_CLR1_g40816 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_809, A2 => hcountintern(6), B1 => TL01_CLR1_n_1014, B2 => TL01_CLR1_n_82, ZN => TL01_CLR1_n_1187);
  TL01_CLR1_g40817 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_990, A2 => TL01_CLR1_n_823, B1 => TL01_CLR1_n_1006, B2 => TL01_CLR1_n_756, C1 => TL01_CLR1_n_43, C2 => TL01_CLR1_n_492, ZN => TL01_CLR1_n_1186);
  TL01_CLR1_g40818 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_1035, A2 => TL01_CLR1_n_739, B => TL01_CLR1_n_1118, ZN => TL01_CLR1_n_1185);
  TL01_CLR1_g40819 : OA22D0BWP7T port map(A1 => TL01_CLR1_n_1107, A2 => TL01_CLR1_n_876, B1 => TL01_CLR1_n_680, B2 => TL01_CLR1_n_830, Z => TL01_CLR1_n_1184);
  TL01_CLR1_g40820 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_910, A2 => TL01_CLR1_n_905, B1 => TL01_CLR1_n_1102, B2 => TL01_CLR1_n_681, ZN => TL01_CLR1_n_1183);
  TL01_CLR1_g40821 : IOA21D1BWP7T port map(A1 => TL01_CLR1_n_1045, A2 => TL01_CLR1_n_82, B => TL01_CLR1_n_1083, ZN => TL01_CLR1_n_1182);
  TL01_CLR1_g40822 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_1108, A2 => TL01_CLR1_n_1076, B1 => TL01_CLR1_n_962, B2 => TL01_CLR1_n_830, ZN => TL01_CLR1_n_1181);
  TL01_CLR1_g40823 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_754, A2 => TL01_CLR1_n_233, B1 => TL01_CLR1_n_1079, B2 => TL01_CLR1_n_379, ZN => TL01_CLR1_n_1180);
  TL01_CLR1_g40824 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_1079, A2 => TL01_CLR1_n_232, B1 => TL01_CLR1_n_754, B2 => TL01_CLR1_n_368, ZN => TL01_CLR1_n_1179);
  TL01_CLR1_g40825 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1105, A2 => TL01_CLR1_n_820, B1 => TL01_CLR1_n_1075, B2 => TL01_CLR1_n_600, ZN => TL01_CLR1_n_1178);
  TL01_CLR1_g40826 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1103, A2 => TL01_CLR1_n_813, B1 => TL01_CLR1_n_972, B2 => TL01_CLR1_n_680, ZN => TL01_CLR1_n_1177);
  TL01_CLR1_g40827 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_1095, A2 => TL01_CLR1_n_819, B1 => TL01_CLR1_n_1036, B2 => TL01_CLR1_n_658, ZN => TL01_CLR1_n_1176);
  TL01_CLR1_g40828 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1089, A2 => TL01_CLR1_n_1093, B1 => TL01_CLR1_n_1100, B2 => TL01_CLR1_n_675, ZN => TL01_CLR1_n_1175);
  TL01_CLR1_g40829 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_1078, A2 => TL01_CLR1_n_235, B1 => TL01_CLR1_n_754, B2 => TL01_CLR1_n_745, ZN => TL01_CLR1_n_1174);
  TL01_CLR1_g40830 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_1079, A2 => TL01_CLR1_n_377, B1 => TL01_CLR1_n_753, B2 => TL01_CLR1_n_234, ZN => TL01_CLR1_n_1173);
  TL01_CLR1_g40831 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_971, A2 => char1posy(7), B1 => TL01_CLR1_n_971, B2 => char1posy(7), ZN => TL01_CLR1_n_1200);
  TL01_CLR1_g40832 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_968, A2 => char2posx(7), B1 => TL01_CLR1_n_968, B2 => char2posx(7), ZN => TL01_CLR1_n_1199);
  TL01_CLR1_g40833 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_973, A2 => char1posx(7), B1 => TL01_CLR1_n_973, B2 => char1posx(7), ZN => TL01_CLR1_n_1198);
  TL01_CLR1_g40834 : NR3D0BWP7T port map(A1 => TL01_CLR1_n_1081, A2 => TL01_CLR1_n_812, A3 => TL01_CLR1_n_484, ZN => TL01_CLR1_n_1197);
  TL01_CLR1_g40835 : NR3D0BWP7T port map(A1 => TL01_CLR1_n_1081, A2 => TL01_CLR1_n_740, A3 => TL01_CLR1_n_682, ZN => TL01_CLR1_n_1195);
  TL01_CLR1_g40836 : INVD1BWP7T port map(I => TL01_CLR1_n_1159, ZN => TL01_CLR1_n_1160);
  TL01_CLR1_g40837 : INVD0BWP7T port map(I => TL01_CLR1_n_1157, ZN => TL01_CLR1_n_1156);
  TL01_CLR1_g40838 : INVD0BWP7T port map(I => TL01_CLR1_n_1155, ZN => TL01_CLR1_n_1154);
  TL01_CLR1_g40839 : INVD0BWP7T port map(I => TL01_CLR1_n_1153, ZN => TL01_CLR1_n_1152);
  TL01_CLR1_g40840 : INVD0BWP7T port map(I => TL01_CLR1_n_1151, ZN => TL01_CLR1_n_1150);
  TL01_CLR1_g40841 : HA1D0BWP7T port map(A => TL01_CLR1_n_74, B => TL01_CLR1_n_835, CO => TL01_CLR1_n_1148, S => TL01_CLR1_n_1172);
  TL01_CLR1_g40842 : HA1D0BWP7T port map(A => TL01_CLR1_n_98, B => TL01_CLR1_n_833, CO => TL01_CLR1_n_1147, S => TL01_CLR1_n_1171);
  TL01_CLR1_g40843 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_564, A2 => TL01_CLR1_n_407, B1 => TL01_CLR1_n_484, B2 => TL01_CLR1_n_321, C => TL01_CLR1_n_1064, ZN => TL01_CLR1_n_1146);
  TL01_CLR1_g40844 : AO211D0BWP7T port map(A1 => TL01_CLR1_n_717, A2 => TL01_CLR1_n_602, B => TL01_CLR1_n_1002, C => TL01_CLR1_n_825, Z => TL01_CLR1_n_1145);
  TL01_CLR1_g40845 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_812, A2 => TL01_CLR1_n_547, B1 => TL01_CLR1_n_484, B2 => TL01_CLR1_n_286, C => TL01_CLR1_n_1065, ZN => TL01_CLR1_n_1144);
  TL01_CLR1_g40846 : IAO21D0BWP7T port map(A1 => TL01_CLR1_n_985, A2 => TL01_CLR1_n_825, B => TL01_CLR1_n_1036, ZN => TL01_CLR1_n_1143);
  TL01_CLR1_g40847 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_724, A2 => TL01_CLR1_n_288, B1 => TL01_CLR1_n_485, B2 => TL01_CLR1_n_283, C => TL01_CLR1_n_1067, ZN => TL01_CLR1_n_1142);
  TL01_CLR1_g40848 : CKAN2D1BWP7T port map(A1 => TL01_CLR1_n_1012, A2 => TL01_CLR1_n_154, Z => TL01_CLR1_n_1141);
  TL01_CLR1_g40849 : INR2XD0BWP7T port map(A1 => TL01_CLR1_n_981, B1 => char2posy(7), ZN => TL01_CLR1_n_1170);
  TL01_CLR1_g40850 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_973, B1 => char1posx(7), ZN => TL01_CLR1_n_1169);
  TL01_CLR1_g40851 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_955, A2 => TL01_CLR1_n_326, B1 => TL01_CLR1_n_618, B2 => TL01_CLR1_n_433, C => TL01_CLR1_n_560, ZN => TL01_CLR1_n_1168);
  TL01_CLR1_g40852 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_971, B1 => char1posy(7), ZN => TL01_CLR1_n_1167);
  TL01_CLR1_g40853 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_968, B1 => char2posx(7), ZN => TL01_CLR1_n_1166);
  TL01_CLR1_g40854 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_1016, A2 => TL01_CLR1_n_59, ZN => TL01_CLR1_n_1165);
  TL01_CLR1_g40855 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1015, A2 => vcountintern(7), ZN => TL01_CLR1_n_1164);
  TL01_CLR1_g40857 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_981, B1 => char2posy(7), ZN => TL01_CLR1_n_1163);
  TL01_CLR1_g40858 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_1113, A2 => TL01_CLR1_n_800, ZN => TL01_CLR1_n_1162);
  TL01_CLR1_g40859 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1111, A2 => TL01_CLR1_n_800, ZN => TL01_CLR1_n_1161);
  TL01_CLR1_g40860 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1110, A2 => TL01_CLR1_n_800, ZN => TL01_CLR1_n_1159);
  TL01_CLR1_g40861 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_1091, A2 => TL01_CLR1_n_493, ZN => TL01_CLR1_n_1158);
  TL01_CLR1_g40862 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_1113, A2 => TL01_CLR1_n_801, ZN => TL01_CLR1_n_1157);
  TL01_CLR1_g40863 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1111, A2 => TL01_CLR1_n_801, ZN => TL01_CLR1_n_1155);
  TL01_CLR1_g40864 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1087, A2 => TL01_CLR1_n_562, ZN => TL01_CLR1_n_1153);
  TL01_CLR1_g40865 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_1112, A2 => TL01_CLR1_n_800, ZN => TL01_CLR1_n_1151);
  TL01_CLR1_g40866 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_1112, A2 => TL01_CLR1_n_801, ZN => TL01_CLR1_n_1149);
  TL01_CLR1_g40867 : NR4D0BWP7T port map(A1 => TL01_CLR1_n_852, A2 => TL01_CLR1_n_927, A3 => TL01_CLR1_n_778, A4 => TL01_CLR1_n_765, ZN => TL01_CLR1_n_1139);
  TL01_CLR1_g40868 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_478, A2 => TL01_CLR1_n_368, B => TL01_CLR1_n_1105, ZN => TL01_CLR1_n_1138);
  TL01_CLR1_g40869 : IND4D0BWP7T port map(A1 => TL01_CLR1_n_692, B1 => TL01_CLR1_n_806, B2 => TL01_CLR1_n_976, B3 => TL01_CLR1_n_1013, ZN => TL01_CLR1_n_1137);
  TL01_CLR1_g40870 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_964, A2 => TL01_CLR1_n_966, B => TL01_CLR1_n_1090, ZN => TL01_CLR1_n_1136);
  TL01_CLR1_g40871 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_964, A2 => char2perc(0), B => TL01_CLR1_n_1090, ZN => TL01_CLR1_n_1135);
  TL01_CLR1_g40872 : AOI211XD0BWP7T port map(A1 => TL01_CLR1_n_799, A2 => TL01_CLR1_n_408, B => TL01_CLR1_n_987, C => TL01_CLR1_n_700, ZN => TL01_CLR1_n_1134);
  TL01_CLR1_g40873 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_912, A2 => char1perc(0), B => TL01_CLR1_n_1090, ZN => TL01_CLR1_n_1133);
  TL01_CLR1_g40874 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_738, A2 => TL01_CLR1_n_326, B1 => TL01_CLR1_n_996, B2 => TL01_CLR1_n_560, ZN => TL01_CLR1_n_1132);
  TL01_CLR1_g40875 : OA21D0BWP7T port map(A1 => TL01_CLR1_n_972, A2 => TL01_CLR1_n_674, B => TL01_CLR1_n_1103, Z => TL01_CLR1_n_1131);
  TL01_CLR1_g40876 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_698, A2 => TL01_CLR1_n_593, B => TL01_CLR1_n_1100, ZN => TL01_CLR1_n_1130);
  TL01_CLR1_g40877 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_994, A2 => TL01_CLR1_n_752, A3 => TL01_CLR1_n_283, ZN => TL01_CLR1_n_1129);
  TL01_CLR1_g40878 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_1036, A2 => TL01_CLR1_n_600, B1 => TL01_CLR1_n_1042, B2 => TL01_CLR1_n_620, ZN => TL01_CLR1_n_1128);
  TL01_CLR1_g40879 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_900, A2 => TL01_CLR1_n_963, B => TL01_CLR1_n_1089, ZN => TL01_CLR1_n_1127);
  TL01_CLR1_g40880 : OA21D0BWP7T port map(A1 => TL01_CLR1_n_803, A2 => TL01_CLR1_n_106, B => TL01_CLR1_n_1015, Z => TL01_CLR1_n_1126);
  TL01_CLR1_g40881 : OAI31D0BWP7T port map(A1 => TL01_CLR1_n_764, A2 => TL01_CLR1_n_774, A3 => TL01_CLR1_n_932, B => TL01_CLR1_n_492, ZN => TL01_CLR1_n_1125);
  TL01_CLR1_g40882 : OAI32D1BWP7T port map(A1 => orientationp1, A2 => TL01_CLR1_char1_sprite_sprite_0, A3 => TL01_CLR1_n_936, B1 => TL01_CLR1_n_1010, B2 => TL01_CLR1_n_1018, ZN => TL01_CLR1_n_1124);
  TL01_CLR1_g40883 : MAOI222D1BWP7T port map(A => TL01_CLR1_n_1004, B => TL01_CLR1_n_610, C => hcountintern(5), ZN => TL01_CLR1_n_1123);
  TL01_CLR1_g40884 : OA221D0BWP7T port map(A1 => TL01_CLR1_n_1032, A2 => TL01_CLR1_n_238, B1 => TL01_CLR1_n_235, B2 => TL01_CLR1_n_811, C => TL01_CLR1_n_787, Z => TL01_CLR1_n_1122);
  TL01_CLR1_g40885 : AO221D0BWP7T port map(A1 => TL01_CLR1_n_952, A2 => TL01_CLR1_n_620, B1 => TL01_CLR1_n_775, B2 => TL01_CLR1_n_751, C => TL01_CLR1_n_992, Z => TL01_CLR1_n_1121);
  TL01_CLR1_g40886 : AOI211XD0BWP7T port map(A1 => TL01_CLR1_n_675, A2 => TL01_CLR1_n_310, B => TL01_CLR1_n_1000, C => TL01_CLR1_n_868, ZN => TL01_CLR1_n_1120);
  TL01_CLR1_g40887 : AO221D0BWP7T port map(A1 => TL01_CLR1_n_1010, A2 => TL01_CLR1_n_576, B1 => TL01_CLR1_n_575, B2 => TL01_CLR1_n_911, C => TL01_CLR1_n_810, Z => TL01_CLR1_n_1119);
  TL01_CLR1_g40888 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_977, A2 => TL01_CLR1_n_675, B1 => TL01_CLR1_n_1041, B2 => TL01_CLR1_n_822, ZN => TL01_CLR1_n_1118);
  TL01_CLR1_g40889 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_977, A2 => TL01_CLR1_n_681, B1 => TL01_CLR1_n_1041, B2 => TL01_CLR1_n_878, ZN => TL01_CLR1_n_1117);
  TL01_CLR1_g40890 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_999, A2 => TL01_CLR1_n_59, B1 => TL01_CLR1_n_607, B2 => TL01_CLR1_n_528, ZN => TL01_CLR1_n_1140);
  TL01_CLR1_g40892 : INVD0BWP7T port map(I => TL01_CLR1_n_1100, ZN => TL01_CLR1_n_1099);
  TL01_CLR1_g40893 : INVD0BWP7T port map(I => TL01_CLR1_n_1098, ZN => TL01_CLR1_n_1097);
  TL01_CLR1_g40894 : INVD1BWP7T port map(I => TL01_CLR1_n_1096, ZN => TL01_CLR1_n_1095);
  TL01_CLR1_g40895 : INVD0BWP7T port map(I => TL01_CLR1_n_1094, ZN => TL01_CLR1_n_1093);
  TL01_CLR1_g40896 : INVD0BWP7T port map(I => TL01_CLR1_n_1092, ZN => TL01_CLR1_n_1091);
  TL01_CLR1_g40897 : INVD1BWP7T port map(I => TL01_CLR1_n_1090, ZN => TL01_CLR1_n_1089);
  TL01_CLR1_g40898 : INVD0BWP7T port map(I => TL01_CLR1_n_1088, ZN => TL01_CLR1_n_1087);
  TL01_CLR1_g40899 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1011, A2 => TL01_CLR1_n_827, ZN => TL01_CLR1_n_1086);
  TL01_CLR1_g40900 : OA221D0BWP7T port map(A1 => TL01_CLR1_n_50, A2 => TL01_CLR1_n_911, B1 => TL01_CLR1_n_72, B2 => TL01_CLR1_char1_sprite_sprite_0, C => TL01_CLR1_n_1009, Z => TL01_CLR1_n_1085);
  TL01_CLR1_g40901 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1009, A2 => TL01_CLR1_n_911, ZN => TL01_CLR1_n_1084);
  TL01_CLR1_g40902 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_1039, A2 => TL01_CLR1_n_975, ZN => TL01_CLR1_n_1116);
  TL01_CLR1_g40903 : NR2D0BWP7T port map(A1 => TL01_CLR1_n_1032, A2 => TL01_CLR1_n_373, ZN => TL01_CLR1_n_1115);
  TL01_CLR1_g40904 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_46, A2 => char2perc(0), ZN => TL01_CLR1_n_1114);
  TL01_CLR1_g40905 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1051, A2 => TL01_CLR1_n_632, ZN => TL01_CLR1_n_1113);
  TL01_CLR1_g40906 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1051, A2 => TL01_CLR1_n_631, ZN => TL01_CLR1_n_1112);
  TL01_CLR1_g40907 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_1046, A2 => TL01_CLR1_n_631, ZN => TL01_CLR1_n_1111);
  TL01_CLR1_g40908 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_1046, A2 => TL01_CLR1_n_632, ZN => TL01_CLR1_n_1110);
  TL01_CLR1_g40909 : INR2XD0BWP7T port map(A1 => TL01_CLR1_n_661, B1 => TL01_CLR1_n_1010, ZN => TL01_CLR1_n_1109);
  TL01_CLR1_g40910 : INR2D1BWP7T port map(A1 => TL01_CLR1_n_1047, B1 => char2perc(0), ZN => TL01_CLR1_n_1108);
  TL01_CLR1_g40911 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_1048, B1 => char2perc(0), ZN => TL01_CLR1_n_1107);
  TL01_CLR1_g40912 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1050, A2 => char2perc(0), ZN => TL01_CLR1_n_1106);
  TL01_CLR1_g40913 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1052, A2 => TL01_CLR1_n_960, ZN => TL01_CLR1_n_1105);
  TL01_CLR1_g40914 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1032, A2 => TL01_CLR1_n_820, ZN => TL01_CLR1_n_1104);
  TL01_CLR1_g40915 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1052, A2 => TL01_CLR1_n_959, ZN => TL01_CLR1_n_1103);
  TL01_CLR1_g40916 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_1049, A2 => TL01_CLR1_n_959, ZN => TL01_CLR1_n_1102);
  TL01_CLR1_g40917 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1050, A2 => FE_DBTN4_char2perc_0, ZN => TL01_CLR1_n_1101);
  TL01_CLR1_g40918 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_1048, A2 => char2perc(0), ZN => TL01_CLR1_n_1100);
  TL01_CLR1_g40919 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_1049, A2 => TL01_CLR1_n_960, ZN => TL01_CLR1_n_1098);
  TL01_CLR1_g40920 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1031, A2 => TL01_CLR1_n_565, ZN => TL01_CLR1_n_1096);
  TL01_CLR1_g40921 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1047, A2 => char2perc(0), ZN => TL01_CLR1_n_1094);
  TL01_CLR1_g40922 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_1039, A2 => TL01_CLR1_n_974, ZN => TL01_CLR1_n_1092);
  TL01_CLR1_g40923 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_1033, A2 => TL01_CLR1_n_846, ZN => TL01_CLR1_n_1090);
  TL01_CLR1_g40924 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_46, A2 => FE_DBTN4_char2perc_0, ZN => TL01_CLR1_n_1088);
  TL01_CLR1_g40925 : INVD0BWP7T port map(I => TL01_CLR1_n_1079, ZN => TL01_CLR1_n_1078);
  TL01_CLR1_g40926 : INVD0BWP7T port map(I => TL01_CLR1_n_1076, ZN => TL01_CLR1_n_1077);
  TL01_CLR1_g40927 : INVD0BWP7T port map(I => TL01_CLR1_n_45, ZN => TL01_CLR1_n_1075);
  TL01_CLR1_g40928 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_508, A2 => TL01_CLR1_n_813, B => TL01_CLR1_n_921, C => TL01_CLR1_n_940, ZN => TL01_CLR1_n_1074);
  TL01_CLR1_g40929 : OAI31D0BWP7T port map(A1 => TL01_CLR1_n_776, A2 => TL01_CLR1_n_933, A3 => TL01_CLR1_n_895, B => TL01_CLR1_n_410, ZN => TL01_CLR1_n_1073);
  TL01_CLR1_g40930 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_906, A2 => TL01_CLR1_n_315, B1 => TL01_CLR1_n_838, B2 => TL01_CLR1_n_310, C => TL01_CLR1_n_882, ZN => TL01_CLR1_n_1072);
  TL01_CLR1_g40931 : ND4D0BWP7T port map(A1 => TL01_CLR1_n_1009, A2 => TL01_CLR1_n_725, A3 => TL01_CLR1_char1_sprite_sprite_1, A4 => orientationp1, ZN => TL01_CLR1_n_1071);
  TL01_CLR1_g40932 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_455, A2 => TL01_CLR1_n_519, B => TL01_CLR1_n_1010, ZN => TL01_CLR1_n_1070);
  TL01_CLR1_g40933 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_558, A2 => TL01_CLR1_n_368, B1 => TL01_CLR1_n_314, B2 => TL01_CLR1_n_559, C => TL01_CLR1_n_1025, ZN => TL01_CLR1_n_1069);
  TL01_CLR1_g40934 : AOI31D0BWP7T port map(A1 => TL01_CLR1_n_745, A2 => TL01_CLR1_n_511, A3 => TL01_CLR1_n_306, B => TL01_CLR1_n_1040, ZN => TL01_CLR1_n_1068);
  TL01_CLR1_g40935 : AOI211XD0BWP7T port map(A1 => TL01_CLR1_n_906, A2 => TL01_CLR1_n_307, B => TL01_CLR1_n_793, C => TL01_CLR1_n_707, ZN => TL01_CLR1_n_1067);
  TL01_CLR1_g40936 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_942, A2 => TL01_CLR1_n_740, B1 => TL01_CLR1_n_812, B2 => TL01_CLR1_n_379, ZN => TL01_CLR1_n_1066);
  TL01_CLR1_g40937 : OAI222D0BWP7T port map(A1 => TL01_CLR1_n_965, A2 => TL01_CLR1_n_238, B1 => TL01_CLR1_n_402, B2 => TL01_CLR1_n_718, C1 => TL01_CLR1_n_311, C2 => TL01_CLR1_n_559, ZN => TL01_CLR1_n_1065);
  TL01_CLR1_g40938 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_724, A2 => TL01_CLR1_n_398, B1 => TL01_CLR1_n_413, B2 => TL01_CLR1_n_907, C => TL01_CLR1_n_650, ZN => TL01_CLR1_n_1064);
  TL01_CLR1_g40939 : AOI31D0BWP7T port map(A1 => TL01_CLR1_n_694, A2 => TL01_CLR1_n_283, A3 => TL01_CLR1_n_375, B => TL01_CLR1_n_1043, ZN => TL01_CLR1_n_1063);
  TL01_CLR1_g40940 : AOI31D0BWP7T port map(A1 => TL01_CLR1_n_883, A2 => TL01_CLR1_n_752, A3 => TL01_CLR1_n_283, B => TL01_CLR1_n_896, ZN => TL01_CLR1_n_1062);
  TL01_CLR1_g40941 : OAI31D0BWP7T port map(A1 => orientationp2, A2 => TL01_CLR1_char2_sprite_sprite_0, A3 => TL01_CLR1_n_848, B => TL01_CLR1_n_1017, ZN => TL01_CLR1_n_1061);
  TL01_CLR1_g40942 : AOI31D0BWP7T port map(A1 => TL01_CLR1_n_849, A2 => TL01_CLR1_n_518, A3 => TL01_CLR1_char1_sprite_sprite_1, B => TL01_CLR1_n_1010, ZN => TL01_CLR1_n_1060);
  TL01_CLR1_g40943 : AOI31D0BWP7T port map(A1 => TL01_CLR1_n_662, A2 => TL01_CLR1_n_566, A3 => TL01_CLR1_n_71, B => TL01_CLR1_n_1021, ZN => TL01_CLR1_n_1059);
  TL01_CLR1_g40944 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_906, A2 => TL01_CLR1_n_312, B1 => TL01_CLR1_n_624, B2 => TL01_CLR1_n_734, C1 => TL01_CLR1_n_763, C2 => TL01_CLR1_n_194, ZN => TL01_CLR1_n_1058);
  TL01_CLR1_g40945 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_376, A2 => TL01_CLR1_n_811, B => TL01_CLR1_n_988, C => TL01_CLR1_n_847, ZN => TL01_CLR1_n_1057);
  TL01_CLR1_g40946 : OAI33D1BWP7T port map(A1 => TL01_CLR1_n_400, A2 => TL01_CLR1_n_394, A3 => TL01_CLR1_n_899, B1 => TL01_CLR1_n_409, B2 => TL01_CLR1_n_547, B3 => TL01_CLR1_n_739, ZN => TL01_CLR1_n_1056);
  TL01_CLR1_g40947 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_824, A2 => char2posx(6), B1 => TL01_CLR1_n_824, B2 => char2posx(6), ZN => TL01_CLR1_n_1083);
  TL01_CLR1_g40948 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_826, A2 => char1posx(6), B1 => TL01_CLR1_n_826, B2 => char1posx(6), ZN => TL01_CLR1_n_1082);
  TL01_CLR1_g40949 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_965, A2 => TL01_CLR1_n_962, A3 => TL01_CLR1_n_621, ZN => TL01_CLR1_n_1081);
  TL01_CLR1_g40950 : IND3D1BWP7T port map(A1 => TL01_CLR1_n_974, B1 => TL01_CLR1_n_729, B2 => TL01_CLR1_n_960, ZN => TL01_CLR1_n_1080);
  TL01_CLR1_g40951 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_965, A2 => TL01_CLR1_n_721, A3 => TL01_CLR1_n_621, ZN => TL01_CLR1_n_1079);
  TL01_CLR1_g40952 : IND4D0BWP7T port map(A1 => TL01_CLR1_n_752, B1 => TL01_CLR1_n_561, B2 => TL01_CLR1_n_626, B3 => TL01_CLR1_n_922, ZN => TL01_CLR1_n_1076);
  TL01_CLR1_g40954 : CKND1BWP7T port map(I => TL01_CLR1_n_1044, ZN => TL01_CLR1_n_1043);
  TL01_CLR1_g40955 : INVD0BWP7T port map(I => TL01_CLR1_n_1034, ZN => TL01_CLR1_n_1035);
  TL01_CLR1_g40956 : INVD1BWP7T port map(I => TL01_CLR1_n_1033, ZN => TL01_CLR1_n_1032);
  TL01_CLR1_g40957 : INVD0BWP7T port map(I => TL01_CLR1_n_1031, ZN => TL01_CLR1_n_1030);
  TL01_CLR1_g40958 : INVD0BWP7T port map(I => TL01_CLR1_n_1029, ZN => TL01_CLR1_n_1028);
  TL01_CLR1_g40959 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_913, A2 => vcountintern(7), Z => TL01_CLR1_n_1027);
  TL01_CLR1_g40960 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_724, A2 => TL01_CLR1_n_405, B1 => TL01_CLR1_n_413, B2 => TL01_CLR1_n_621, C => TL01_CLR1_n_935, ZN => TL01_CLR1_n_1026);
  TL01_CLR1_g40961 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_812, A2 => TL01_CLR1_n_629, B1 => TL01_CLR1_n_484, B2 => TL01_CLR1_n_310, C => TL01_CLR1_n_779, ZN => TL01_CLR1_n_1025);
  TL01_CLR1_g40962 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_198, A2 => TL01_CLR1_n_679, B => TL01_CLR1_n_875, C => TL01_CLR1_n_767, ZN => TL01_CLR1_n_1024);
  TL01_CLR1_g40963 : AOI31D0BWP7T port map(A1 => TL01_CLR1_n_784, A2 => TL01_CLR1_n_623, A3 => TL01_CLR1_n_600, B => TL01_CLR1_n_781, ZN => TL01_CLR1_n_1023);
  TL01_CLR1_g40964 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_886, A2 => TL01_CLR1_n_945, ZN => TL01_CLR1_n_1022);
  TL01_CLR1_g40965 : NR2D0BWP7T port map(A1 => TL01_CLR1_char2_sprite_sprite_0, A2 => TL01_CLR1_n_970, ZN => TL01_CLR1_n_1021);
  TL01_CLR1_g40966 : AN2D0BWP7T port map(A1 => TL01_CLR1_n_914, A2 => TL01_CLR1_n_169, Z => TL01_CLR1_n_1020);
  TL01_CLR1_g40967 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_980, A2 => TL01_CLR1_n_603, Z => TL01_CLR1_n_1019);
  TL01_CLR1_g40969 : INR2XD0BWP7T port map(A1 => char2posx(6), B1 => TL01_CLR1_n_824, ZN => TL01_CLR1_n_1055);
  TL01_CLR1_g40970 : INR2XD0BWP7T port map(A1 => char1posx(6), B1 => TL01_CLR1_n_826, ZN => TL01_CLR1_n_1054);
  TL01_CLR1_g40971 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_920, A2 => TL01_CLR1_n_154, ZN => TL01_CLR1_n_1053);
  TL01_CLR1_g40972 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_975, A2 => TL01_CLR1_n_729, ZN => TL01_CLR1_n_1052);
  TL01_CLR1_g40973 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_966, A2 => TL01_CLR1_n_727, ZN => TL01_CLR1_n_1051);
  TL01_CLR1_g40974 : INR2D1BWP7T port map(A1 => TL01_CLR1_n_757, B1 => TL01_CLR1_n_967, ZN => TL01_CLR1_n_1050);
  TL01_CLR1_g40975 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_974, A2 => TL01_CLR1_n_729, Z => TL01_CLR1_n_1049);
  TL01_CLR1_g40976 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_967, A2 => TL01_CLR1_n_757, ZN => TL01_CLR1_n_1048);
  TL01_CLR1_g40977 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_967, A2 => TL01_CLR1_n_757, ZN => TL01_CLR1_n_1047);
  TL01_CLR1_g40978 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_966, A2 => TL01_CLR1_n_726, ZN => TL01_CLR1_n_1046);
  TL01_CLR1_g40979 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_917, A2 => TL01_CLR1_n_154, ZN => TL01_CLR1_n_1045);
  TL01_CLR1_g40980 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_900, A2 => TL01_CLR1_n_950, ZN => TL01_CLR1_n_1044);
  TL01_CLR1_g40981 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_901, A2 => TL01_CLR1_n_979, ZN => TL01_CLR1_n_1042);
  TL01_CLR1_g40982 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_901, A2 => TL01_CLR1_n_983, ZN => TL01_CLR1_n_1041);
  TL01_CLR1_g40983 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_901, A2 => TL01_CLR1_n_978, ZN => TL01_CLR1_n_1040);
  TL01_CLR1_g40984 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_959, A2 => TL01_CLR1_n_729, ZN => TL01_CLR1_n_1039);
  TL01_CLR1_g40985 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_966, A2 => TL01_CLR1_n_727, ZN => TL01_CLR1_n_1038);
  TL01_CLR1_g40986 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_900, A2 => TL01_CLR1_n_978, ZN => TL01_CLR1_n_1037);
  TL01_CLR1_g40987 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_900, A2 => TL01_CLR1_n_983, ZN => TL01_CLR1_n_1036);
  TL01_CLR1_g40988 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_900, A2 => TL01_CLR1_n_979, ZN => TL01_CLR1_n_1034);
  TL01_CLR1_g40989 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_965, A2 => TL01_CLR1_n_811, ZN => TL01_CLR1_n_1033);
  TL01_CLR1_g40990 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_901, A2 => TL01_CLR1_n_950, ZN => TL01_CLR1_n_1031);
  TL01_CLR1_g40991 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_963, A2 => TL01_CLR1_n_484, ZN => TL01_CLR1_n_1029);
  TL01_CLR1_g40993 : INVD1BWP7T port map(I => TL01_CLR1_n_1010, ZN => TL01_CLR1_n_1009);
  TL01_CLR1_g40994 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_663, A2 => TL01_CLR1_n_872, B1 => TL01_CLR1_n_888, B2 => TL01_CLR1_n_176, ZN => TL01_CLR1_n_1008);
  TL01_CLR1_g40995 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_855, A2 => TL01_CLR1_n_756, B1 => TL01_CLR1_n_823, B2 => TL01_CLR1_n_821, ZN => TL01_CLR1_n_1007);
  TL01_CLR1_g40996 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_402, A2 => TL01_CLR1_n_44, B => TL01_CLR1_n_923, C => TL01_CLR1_n_890, ZN => TL01_CLR1_n_1006);
  TL01_CLR1_g40997 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_814, A2 => TL01_CLR1_n_719, B1 => TL01_CLR1_n_816, B2 => TL01_CLR1_n_287, C1 => TL01_CLR1_n_673, C2 => TL01_CLR1_n_236, ZN => TL01_CLR1_n_1005);
  TL01_CLR1_g40998 : IAO21D0BWP7T port map(A1 => TL01_CLR1_n_696, A2 => hcountintern(4), B => TL01_CLR1_n_938, ZN => TL01_CLR1_n_1004);
  TL01_CLR1_g40999 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_378, A2 => TL01_CLR1_char2_sprite_sprite_1, B => TL01_CLR1_n_969, ZN => TL01_CLR1_n_1003);
  TL01_CLR1_g41000 : NR4D0BWP7T port map(A1 => TL01_CLR1_n_828, A2 => TL01_CLR1_n_602, A3 => TL01_CLR1_n_629, A4 => TL01_CLR1_n_374, ZN => TL01_CLR1_n_1002);
  TL01_CLR1_g41001 : OA221D0BWP7T port map(A1 => TL01_CLR1_n_815, A2 => TL01_CLR1_n_405, B1 => TL01_CLR1_n_309, B2 => TL01_CLR1_n_44, C => TL01_CLR1_n_923, Z => TL01_CLR1_n_1001);
  TL01_CLR1_g41002 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_744, A2 => TL01_CLR1_n_319, B1 => TL01_CLR1_n_313, B2 => TL01_CLR1_n_679, C => TL01_CLR1_n_941, ZN => TL01_CLR1_n_1000);
  TL01_CLR1_g41003 : ND4D0BWP7T port map(A1 => TL01_CLR1_n_785, A2 => TL01_CLR1_n_396, A3 => TL01_CLR1_n_433, A4 => TL01_CLR1_n_148, ZN => TL01_CLR1_n_999);
  TL01_CLR1_g41004 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_744, A2 => TL01_CLR1_n_375, B1 => TL01_CLR1_n_288, B2 => TL01_CLR1_n_798, C => TL01_CLR1_n_858, ZN => TL01_CLR1_n_998);
  TL01_CLR1_g41005 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_716, A2 => TL01_CLR1_n_808, B => TL01_CLR1_n_560, C => TL01_CLR1_n_432, ZN => TL01_CLR1_n_997);
  TL01_CLR1_g41006 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_894, A2 => TL01_CLR1_n_433, B => TL01_CLR1_n_545, ZN => TL01_CLR1_n_996);
  TL01_CLR1_g41007 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_887, A2 => TL01_CLR1_n_840, B => TL01_CLR1_n_42, ZN => TL01_CLR1_n_995);
  TL01_CLR1_g41008 : INR4D0BWP7T port map(A1 => TL01_CLR1_n_690, B1 => TL01_CLR1_n_629, B2 => TL01_CLR1_n_834, B3 => TL01_CLR1_n_602, ZN => TL01_CLR1_n_994);
  TL01_CLR1_g41009 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_816, A2 => TL01_CLR1_n_412, B1 => TL01_CLR1_n_814, B2 => TL01_CLR1_n_489, C1 => TL01_CLR1_n_673, C2 => TL01_CLR1_n_374, ZN => TL01_CLR1_n_993);
  TL01_CLR1_g41010 : AOI31D0BWP7T port map(A1 => TL01_CLR1_n_676, A2 => TL01_CLR1_n_844, A3 => TL01_CLR1_n_581, B => TL01_CLR1_n_818, ZN => TL01_CLR1_n_992);
  TL01_CLR1_g41011 : OA221D0BWP7T port map(A1 => TL01_CLR1_n_813, A2 => TL01_CLR1_n_246, B1 => TL01_CLR1_n_723, B2 => TL01_CLR1_n_44, C => TL01_CLR1_n_921, Z => TL01_CLR1_n_991);
  TL01_CLR1_g41012 : IND4D0BWP7T port map(A1 => TL01_CLR1_n_819, B1 => TL01_CLR1_n_581, B2 => TL01_CLR1_n_907, B3 => TL01_CLR1_n_903, ZN => TL01_CLR1_n_990);
  TL01_CLR1_g41013 : AOI31D0BWP7T port map(A1 => TL01_CLR1_n_842, A2 => TL01_CLR1_n_284, A3 => TL01_CLR1_n_320, B => TL01_CLR1_n_825, ZN => TL01_CLR1_n_989);
  TL01_CLR1_g41014 : ND4D0BWP7T port map(A1 => TL01_CLR1_n_829, A2 => TL01_CLR1_n_745, A3 => TL01_CLR1_n_376, A4 => TL01_CLR1_n_373, ZN => TL01_CLR1_n_988);
  TL01_CLR1_g41015 : AOI32D1BWP7T port map(A1 => TL01_CLR1_n_739, A2 => TL01_CLR1_n_795, A3 => TL01_CLR1_n_687, B1 => TL01_CLR1_n_460, B2 => TL01_CLR1_n_316, ZN => TL01_CLR1_n_987);
  TL01_CLR1_g41016 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_516, A2 => TL01_CLR1_n_925, B1 => TL01_CLR1_char2_sprite_sprite_1, B2 => TL01_CLR1_char2_sprite_sprite_0, ZN => TL01_CLR1_n_986);
  TL01_CLR1_g41017 : OAI32D1BWP7T port map(A1 => TL01_CLR1_n_236, A2 => TL01_CLR1_n_316, A3 => TL01_CLR1_n_841, B1 => TL01_CLR1_n_723, B2 => TL01_CLR1_n_718, ZN => TL01_CLR1_n_985);
  TL01_CLR1_g41018 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_918, A2 => TL01_CLR1_n_725, A3 => TL01_CLR1_n_519, ZN => TL01_CLR1_n_1018);
  TL01_CLR1_g41019 : IAO21D0BWP7T port map(A1 => TL01_CLR1_n_669, A2 => hcountintern(4), B => TL01_CLR1_n_937, ZN => TL01_CLR1_n_984);
  TL01_CLR1_g41020 : IND3D1BWP7T port map(A1 => TL01_CLR1_n_970, B1 => TL01_CLR1_n_566, B2 => TL01_CLR1_n_378, ZN => TL01_CLR1_n_1017);
  TL01_CLR1_g41021 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_759, A2 => char1posy(6), B1 => TL01_CLR1_n_759, B2 => char1posy(6), ZN => TL01_CLR1_n_1016);
  TL01_CLR1_g41022 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_762, A2 => char2posy(6), B1 => TL01_CLR1_n_762, B2 => char2posy(6), ZN => TL01_CLR1_n_1015);
  TL01_CLR1_g41023 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_758, A2 => char1posx(6), B1 => TL01_CLR1_n_758, B2 => char1posx(6), ZN => TL01_CLR1_n_1014);
  TL01_CLR1_g41024 : AOI211XD0BWP7T port map(A1 => TL01_CLR1_n_792, A2 => vcountintern(7), B => TL01_CLR1_n_916, C => TL01_CLR1_n_769, ZN => TL01_CLR1_n_1013);
  TL01_CLR1_g41025 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_761, A2 => char2posx(6), B => TL01_CLR1_n_968, ZN => TL01_CLR1_n_1012);
  TL01_CLR1_g41026 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_884, A2 => vcountintern(4), B1 => TL01_CLR1_n_884, B2 => vcountintern(4), ZN => TL01_CLR1_n_1011);
  TL01_CLR1_g41027 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_885, A2 => vcountintern(4), B1 => TL01_CLR1_n_885, B2 => vcountintern(4), ZN => TL01_CLR1_n_1010);
  TL01_CLR1_g41028 : INVD0BWP7T port map(I => TL01_CLR1_n_970, ZN => TL01_CLR1_n_969);
  TL01_CLR1_g41030 : INVD0BWP7T port map(I => TL01_CLR1_n_963, ZN => TL01_CLR1_n_964);
  TL01_CLR1_g41031 : INVD1BWP7T port map(I => TL01_CLR1_n_961, ZN => TL01_CLR1_n_962);
  TL01_CLR1_g41032 : INVD1BWP7T port map(I => TL01_CLR1_n_960, ZN => TL01_CLR1_n_959);
  TL01_CLR1_g41033 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_804, A2 => TL01_CLR1_n_59, Z => TL01_CLR1_n_958);
  TL01_CLR1_g41034 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_744, A2 => TL01_CLR1_n_402, B1 => TL01_CLR1_n_401, B2 => TL01_CLR1_n_623, C => TL01_CLR1_n_839, ZN => TL01_CLR1_n_957);
  TL01_CLR1_g41035 : AO221D0BWP7T port map(A1 => TL01_CLR1_n_770, A2 => TL01_CLR1_n_491, B1 => TL01_CLR1_n_749, B2 => TL01_CLR1_n_494, C => TL01_CLR1_n_764, Z => TL01_CLR1_n_956);
  TL01_CLR1_g41036 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_834, A2 => TL01_CLR1_n_539, B => TL01_CLR1_n_429, ZN => TL01_CLR1_n_955);
  TL01_CLR1_g41037 : ND2D0BWP7T port map(A1 => TL01_CLR1_n_919, A2 => TL01_CLR1_n_561, ZN => TL01_CLR1_n_954);
  TL01_CLR1_g41038 : IND2D0BWP7T port map(A1 => TL01_CLR1_n_624, B1 => TL01_CLR1_n_908, ZN => TL01_CLR1_n_953);
  TL01_CLR1_g41039 : INR2D1BWP7T port map(A1 => TL01_CLR1_n_630, B1 => TL01_CLR1_n_909, ZN => TL01_CLR1_n_983);
  TL01_CLR1_g41040 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_803, A2 => vcountintern(6), ZN => TL01_CLR1_n_982);
  TL01_CLR1_g41041 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_762, A2 => TL01_CLR1_n_98, Z => TL01_CLR1_n_981);
  TL01_CLR1_g41042 : INR2D1BWP7T port map(A1 => vcountintern(6), B1 => TL01_CLR1_n_804, ZN => TL01_CLR1_n_980);
  TL01_CLR1_g41043 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_630, B1 => TL01_CLR1_n_909, ZN => TL01_CLR1_n_979);
  TL01_CLR1_g41044 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_909, A2 => TL01_CLR1_n_630, ZN => TL01_CLR1_n_978);
  TL01_CLR1_g41045 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_900, A2 => TL01_CLR1_n_601, ZN => TL01_CLR1_n_977);
  TL01_CLR1_g41046 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_794, A2 => TL01_CLR1_n_262, A3 => TL01_CLR1_n_90, ZN => TL01_CLR1_n_976);
  TL01_CLR1_g41047 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_905, A2 => char1perc(0), ZN => TL01_CLR1_n_975);
  TL01_CLR1_g41048 : IND2D1BWP7T port map(A1 => char1perc(0), B1 => TL01_CLR1_n_905, ZN => TL01_CLR1_n_974);
  TL01_CLR1_g41049 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_758, B1 => char1posx(6), ZN => TL01_CLR1_n_973);
  TL01_CLR1_g41050 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_904, A2 => char1perc(0), ZN => TL01_CLR1_n_972);
  TL01_CLR1_g41051 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_759, A2 => TL01_CLR1_n_74, Z => TL01_CLR1_n_971);
  TL01_CLR1_g41052 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_728, A2 => TL01_CLR1_n_516, B => TL01_CLR1_n_71, ZN => TL01_CLR1_n_970);
  TL01_CLR1_g41053 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_761, A2 => char2posx(6), ZN => TL01_CLR1_n_968);
  TL01_CLR1_g41054 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_522, A2 => TL01_CLR1_n_381, B1 => TL01_CLR1_n_422, B2 => TL01_CLR1_n_112, C => TL01_CLR1_n_869, ZN => TL01_CLR1_n_967);
  TL01_CLR1_g41055 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_347, A2 => TL01_CLR1_n_529, B => TL01_CLR1_n_874, C => TL01_CLR1_n_477, ZN => TL01_CLR1_n_966);
  TL01_CLR1_g41056 : CKAN2D1BWP7T port map(A1 => TL01_CLR1_n_908, A2 => TL01_CLR1_n_747, Z => TL01_CLR1_n_965);
  TL01_CLR1_g41057 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_912, A2 => TL01_CLR1_n_623, ZN => TL01_CLR1_n_963);
  TL01_CLR1_g41058 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_912, A2 => TL01_CLR1_n_798, ZN => TL01_CLR1_n_961);
  TL01_CLR1_g41059 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_873, A2 => TL01_CLR1_n_520, A3 => TL01_CLR1_n_454, ZN => TL01_CLR1_n_960);
  TL01_CLR1_g41060 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_368, A2 => TL01_CLR1_n_744, B => TL01_CLR1_n_777, C => TL01_CLR1_n_783, ZN => TL01_CLR1_n_949);
  TL01_CLR1_g41061 : AO21D0BWP7T port map(A1 => TL01_CLR1_n_752, A2 => TL01_CLR1_n_549, B => TL01_CLR1_n_879, Z => TL01_CLR1_n_948);
  TL01_CLR1_g41062 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_811, A2 => TL01_CLR1_n_233, B1 => TL01_CLR1_n_558, B2 => TL01_CLR1_n_309, ZN => TL01_CLR1_n_947);
  TL01_CLR1_g41063 : AOI211XD0BWP7T port map(A1 => TL01_CLR1_n_620, A2 => TL01_CLR1_n_334, B => TL01_CLR1_n_859, C => TL01_CLR1_n_789, ZN => TL01_CLR1_n_946);
  TL01_CLR1_g41064 : ND4D0BWP7T port map(A1 => TL01_CLR1_n_752, A2 => TL01_CLR1_n_309, A3 => TL01_CLR1_n_317, A4 => TL01_CLR1_n_1495, ZN => TL01_CLR1_n_945);
  TL01_CLR1_g41065 : AO31D1BWP7T port map(A1 => TL01_CLR1_n_711, A2 => TL01_CLR1_n_573, A3 => TL01_CLR1_n_545, B => TL01_CLR1_n_626, Z => TL01_CLR1_n_944);
  TL01_CLR1_g41066 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_193, A2 => TL01_CLR1_n_679, B => TL01_CLR1_n_853, C => TL01_CLR1_n_767, ZN => TL01_CLR1_n_943);
  TL01_CLR1_g41067 : NR4D0BWP7T port map(A1 => TL01_CLR1_n_720, A2 => TL01_CLR1_n_722, A3 => TL01_CLR1_n_367, A4 => TL01_CLR1_n_379, ZN => TL01_CLR1_n_942);
  TL01_CLR1_g41068 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_742, A2 => TL01_CLR1_n_285, B1 => TL01_CLR1_n_799, B2 => TL01_CLR1_n_286, ZN => TL01_CLR1_n_941);
  TL01_CLR1_g41069 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_834, A2 => TL01_CLR1_n_512, B => TL01_CLR1_n_673, ZN => TL01_CLR1_n_940);
  TL01_CLR1_g41070 : IOA21D1BWP7T port map(A1 => TL01_CLR1_n_829, A2 => TL01_CLR1_n_572, B => TL01_CLR1_n_836, ZN => TL01_CLR1_n_939);
  TL01_CLR1_g41071 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_705, A2 => TL01_CLR1_n_552, B1 => TL01_CLR1_n_608, B2 => TL01_CLR1_n_596, C1 => TL01_CLR1_n_696, C2 => hcountintern(4), ZN => TL01_CLR1_n_938);
  TL01_CLR1_g41072 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_710, A2 => TL01_CLR1_n_553, B1 => TL01_CLR1_n_609, B2 => TL01_CLR1_n_597, C1 => TL01_CLR1_n_669, C2 => hcountintern(4), ZN => TL01_CLR1_n_937);
  TL01_CLR1_g41073 : AOI32D1BWP7T port map(A1 => TL01_CLR1_n_772, A2 => TL01_CLR1_n_455, A3 => TL01_CLR1_n_519, B1 => TL01_CLR1_n_845, B2 => TL01_CLR1_n_725, ZN => TL01_CLR1_n_936);
  TL01_CLR1_g41074 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_802, A2 => TL01_CLR1_n_399, B1 => TL01_CLR1_n_763, B2 => TL01_CLR1_n_407, C1 => TL01_CLR1_n_580, C2 => TL01_CLR1_n_624, ZN => TL01_CLR1_n_935);
  TL01_CLR1_g41075 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_827, A2 => TL01_CLR1_n_516, B1 => TL01_CLR1_char2_sprite_sprite_1, B2 => orientationp2, ZN => TL01_CLR1_n_934);
  TL01_CLR1_g41076 : OAI32D0BWP7T port map(A1 => TL01_hcount_int(0), A2 => TL01_CLR1_n_561, A3 => TL01_CLR1_n_719, B1 => TL01_CLR1_n_495, B2 => TL01_CLR1_n_676, ZN => TL01_CLR1_n_933);
  TL01_CLR1_g41077 : OAI222D0BWP7T port map(A1 => TL01_CLR1_n_744, A2 => TL01_CLR1_n_486, B1 => TL01_CLR1_n_395, B2 => TL01_CLR1_n_798, C1 => TL01_CLR1_n_401, C2 => TL01_CLR1_n_741, ZN => TL01_CLR1_n_932);
  TL01_CLR1_g41078 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_743, A2 => TL01_CLR1_n_746, B1 => TL01_CLR1_n_742, B2 => TL01_CLR1_n_234, C1 => TL01_CLR1_n_677, C2 => TL01_CLR1_n_412, ZN => TL01_CLR1_n_931);
  TL01_CLR1_g41079 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_644, A2 => TL01_CLR1_n_44, B1 => TL01_CLR1_n_821, B2 => TL01_CLR1_n_488, ZN => TL01_CLR1_n_930);
  TL01_CLR1_g41080 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_802, A2 => TL01_CLR1_n_577, B1 => TL01_CLR1_n_838, B2 => TL01_CLR1_n_286, ZN => TL01_CLR1_n_929);
  TL01_CLR1_g41081 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_309, A2 => TL01_CLR1_n_744, B => TL01_CLR1_n_839, C => TL01_CLR1_n_766, ZN => TL01_CLR1_n_928);
  TL01_CLR1_g41082 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_744, A2 => TL01_CLR1_n_411, B1 => TL01_CLR1_n_798, B2 => TL01_CLR1_n_306, ZN => TL01_CLR1_n_927);
  TL01_CLR1_g41083 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_675, A2 => TL01_CLR1_n_394, B1 => TL01_CLR1_n_799, B2 => TL01_CLR1_n_400, ZN => TL01_CLR1_n_926);
  TL01_CLR1_g41084 : OAI31D0BWP7T port map(A1 => TL01_hcount_int(0), A2 => TL01_CLR1_n_719, A3 => TL01_CLR1_n_750, B => TL01_CLR1_n_818, ZN => TL01_CLR1_n_952);
  TL01_CLR1_g41085 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_846, A2 => TL01_CLR1_n_374, B1 => TL01_CLR1_n_557, B2 => TL01_CLR1_n_236, ZN => TL01_CLR1_n_951);
  TL01_CLR1_g41086 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_909, A2 => TL01_CLR1_n_601, A3 => TL01_CLR1_n_630, ZN => TL01_CLR1_n_950);
  TL01_CLR1_g41087 : INVD0BWP7T port map(I => TL01_CLR1_n_924, ZN => TL01_CLR1_n_925);
  TL01_CLR1_g41088 : INVD1BWP7T port map(I => TL01_CLR1_n_915, ZN => TL01_CLR1_n_916);
  TL01_CLR1_g41089 : INVD1BWP7T port map(I => TL01_CLR1_n_907, ZN => TL01_CLR1_n_906);
  TL01_CLR1_g41090 : INVD0BWP7T port map(I => TL01_CLR1_n_905, ZN => TL01_CLR1_n_904);
  TL01_CLR1_g41091 : INVD0BWP7T port map(I => TL01_CLR1_n_903, ZN => TL01_CLR1_n_902);
  TL01_CLR1_g41092 : INVD1BWP7T port map(I => TL01_CLR1_n_901, ZN => TL01_CLR1_n_900);
  TL01_CLR1_g41093 : IND4D0BWP7T port map(A1 => TL01_CLR1_n_491, B1 => TL01_CLR1_n_495, B2 => TL01_CLR1_n_42, B3 => TL01_CLR1_n_752, ZN => TL01_CLR1_n_899);
  TL01_CLR1_g41096 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_802, B1 => TL01_CLR1_n_686, ZN => TL01_CLR1_n_898);
  TL01_CLR1_g41097 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_742, A2 => TL01_CLR1_n_622, B => TL01_CLR1_n_823, ZN => TL01_CLR1_n_897);
  TL01_CLR1_g41098 : AOI31D0BWP7T port map(A1 => TL01_CLR1_n_385, A2 => TL01_CLR1_n_317, A3 => TL01_CLR1_n_325, B => TL01_CLR1_n_811, ZN => TL01_CLR1_n_896);
  TL01_CLR1_g41099 : AO21D0BWP7T port map(A1 => TL01_CLR1_n_743, A2 => TL01_CLR1_n_488, B => TL01_CLR1_n_843, Z => TL01_CLR1_n_895);
  TL01_CLR1_g41100 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_400, A2 => vcountintern(0), B => TL01_CLR1_n_808, ZN => TL01_CLR1_n_894);
  TL01_CLR1_g41101 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_685, A2 => TL01_CLR1_n_624, B => TL01_CLR1_n_823, ZN => TL01_CLR1_n_893);
  TL01_CLR1_g41102 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_821, A2 => TL01_CLR1_n_749, ZN => TL01_CLR1_n_892);
  TL01_CLR1_g41103 : OA21D0BWP7T port map(A1 => TL01_CLR1_n_458, A2 => TL01_CLR1_n_1494, B => TL01_CLR1_n_791, Z => TL01_CLR1_n_891);
  TL01_CLR1_g41104 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_816, A2 => TL01_CLR1_n_286, ZN => TL01_CLR1_n_890);
  TL01_CLR1_g41106 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_676, A2 => TL01_CLR1_n_403, B1 => TL01_CLR1_n_413, B2 => TL01_CLR1_n_679, C => TL01_CLR1_n_788, ZN => TL01_CLR1_n_889);
  TL01_CLR1_g41107 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_695, A2 => TL01_CLR1_n_611, B1 => TL01_CLR1_n_457, B2 => vcountintern(5), ZN => TL01_CLR1_n_888);
  TL01_CLR1_g41109 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_848, A2 => TL01_CLR1_n_71, ZN => TL01_CLR1_n_924);
  TL01_CLR1_g41110 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_814, A2 => TL01_CLR1_n_283, ZN => TL01_CLR1_n_923);
  TL01_CLR1_g41111 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_799, A2 => TL01_CLR1_n_627, ZN => TL01_CLR1_n_922);
  TL01_CLR1_g41112 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_816, A2 => TL01_CLR1_n_285, ZN => TL01_CLR1_n_921);
  TL01_CLR1_g41113 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_637, A2 => char1posx(5), B => TL01_CLR1_n_826, ZN => TL01_CLR1_n_920);
  TL01_CLR1_g41114 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_821, A2 => TL01_CLR1_n_742, ZN => TL01_CLR1_n_919);
  TL01_CLR1_g41115 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_845, A2 => TL01_CLR1_char1_sprite_sprite_0, ZN => TL01_CLR1_n_918);
  TL01_CLR1_g41116 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_641, A2 => char2posx(5), B => TL01_CLR1_n_824, ZN => TL01_CLR1_n_917);
  TL01_CLR1_g41117 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_796, A2 => FE_OFN3_reset, ZN => TL01_CLR1_n_915);
  TL01_CLR1_g41118 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_635, A2 => char2posy(5), B => TL01_CLR1_n_833, ZN => TL01_CLR1_n_914);
  TL01_CLR1_g41119 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_639, A2 => char1posy(5), B => TL01_CLR1_n_835, ZN => TL01_CLR1_n_913);
  TL01_CLR1_g41120 : CKAN2D1BWP7T port map(A1 => TL01_CLR1_n_844, A2 => TL01_CLR1_n_626, Z => TL01_CLR1_n_912);
  TL01_CLR1_g41121 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_849, A2 => TL01_CLR1_n_519, A3 => TL01_CLR1_n_72, ZN => TL01_CLR1_n_911);
  TL01_CLR1_g41122 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_814, A2 => TL01_CLR1_n_682, ZN => TL01_CLR1_n_910);
  TL01_CLR1_g41123 : AOI211D1BWP7T port map(A1 => TL01_CLR1_n_131, A2 => TL01_CLR1_n_132, B => TL01_CLR1_n_708, C => TL01_CLR1_n_218, ZN => TL01_CLR1_n_909);
  TL01_CLR1_g41124 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_802, A2 => TL01_CLR1_n_564, ZN => TL01_CLR1_n_908);
  TL01_CLR1_g41125 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_802, A2 => TL01_CLR1_n_327, ZN => TL01_CLR1_n_907);
  TL01_CLR1_g41126 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_470, A2 => TL01_CLR1_n_250, B1 => TL01_CLR1_n_506, B2 => TL01_CLR1_n_342, C => TL01_CLR1_n_780, ZN => TL01_CLR1_n_905);
  TL01_CLR1_g41127 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_816, A2 => TL01_CLR1_n_673, ZN => TL01_CLR1_n_903);
  TL01_CLR1_g41128 : OAI221D1BWP7T port map(A1 => TL01_CLR1_n_355, A2 => char1perc(2), B1 => TL01_CLR1_n_191, B2 => TL01_CLR1_n_448, C => TL01_CLR1_n_715, ZN => TL01_CLR1_n_901);
  TL01_CLR1_g41129 : INVD0BWP7T port map(I => TL01_CLR1_n_886, ZN => TL01_CLR1_n_887);
  TL01_CLR1_g41130 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_721, A2 => TL01_CLR1_n_233, B1 => TL01_CLR1_n_564, B2 => TL01_CLR1_n_334, ZN => TL01_CLR1_n_882);
  TL01_CLR1_g41131 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_619, A2 => TL01_CLR1_n_749, B1 => TL01_CLR1_n_679, B2 => TL01_CLR1_n_403, ZN => TL01_CLR1_n_881);
  TL01_CLR1_g41132 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_751, A2 => TL01_CLR1_n_367, B => TL01_CLR1_n_817, ZN => TL01_CLR1_n_880);
  TL01_CLR1_g41133 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_572, A2 => TL01_CLR1_n_238, B => TL01_CLR1_n_811, ZN => TL01_CLR1_n_879);
  TL01_CLR1_g41134 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_557, A2 => TL01_CLR1_n_233, B => TL01_CLR1_n_814, ZN => TL01_CLR1_n_878);
  TL01_CLR1_g41135 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_740, A2 => TL01_CLR1_n_235, B => TL01_CLR1_n_681, ZN => TL01_CLR1_n_877);
  TL01_CLR1_g41136 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_557, A2 => TL01_CLR1_n_376, B => TL01_CLR1_n_814, ZN => TL01_CLR1_n_876);
  TL01_CLR1_g41137 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_743, A2 => TL01_CLR1_n_285, B1 => TL01_CLR1_n_742, B2 => TL01_CLR1_n_286, ZN => TL01_CLR1_n_875);
  TL01_CLR1_g41138 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_652, A2 => char2perc(1), B1 => TL01_CLR1_n_544, B2 => FE_DBTN9_char2perc_5, C1 => TL01_CLR1_n_445, C2 => char2perc(5), ZN => TL01_CLR1_n_874);
  TL01_CLR1_g41139 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_548, A2 => char1perc(7), B1 => TL01_CLR1_n_383, B2 => TL01_CLR1_n_451, C => TL01_CLR1_n_714, ZN => TL01_CLR1_n_873);
  TL01_CLR1_g41140 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_695, A2 => vcountintern(5), B1 => TL01_CLR1_n_457, B2 => vcountintern(4), ZN => TL01_CLR1_n_872);
  TL01_CLR1_g41141 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_666, A2 => vcountintern(5), B1 => TL01_CLR1_n_583, B2 => vcountintern(4), ZN => TL01_CLR1_n_871);
  TL01_CLR1_g41142 : OAI222D0BWP7T port map(A1 => TL01_CLR1_n_720, A2 => TL01_CLR1_n_600, B1 => TL01_CLR1_n_313, B2 => TL01_CLR1_n_559, C1 => TL01_CLR1_n_485, C2 => TL01_CLR1_n_306, ZN => TL01_CLR1_n_870);
  TL01_CLR1_g41143 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_297, A2 => TL01_CLR1_n_346, B1 => TL01_CLR1_n_242, B2 => TL01_CLR1_n_524, C => TL01_CLR1_n_709, ZN => TL01_CLR1_n_869);
  TL01_CLR1_g41144 : OAI222D0BWP7T port map(A1 => TL01_CLR1_n_676, A2 => TL01_CLR1_n_322, B1 => TL01_CLR1_n_193, B2 => TL01_CLR1_n_44, C1 => TL01_CLR1_n_198, C2 => TL01_CLR1_n_561, ZN => TL01_CLR1_n_868);
  TL01_CLR1_g41145 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_665, A2 => hcountintern(5), B1 => TL01_CLR1_n_461, B2 => hcountintern(4), ZN => TL01_CLR1_n_867);
  TL01_CLR1_g41146 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_668, A2 => hcountintern(5), B1 => TL01_CLR1_n_459, B2 => hcountintern(4), ZN => TL01_CLR1_n_866);
  TL01_CLR1_g41147 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_745, A2 => TL01_CLR1_n_558, B1 => TL01_CLR1_n_621, B2 => TL01_CLR1_n_309, ZN => TL01_CLR1_n_865);
  TL01_CLR1_g41148 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_720, A2 => TL01_CLR1_n_620, B1 => TL01_CLR1_n_557, B2 => TL01_CLR1_n_321, ZN => TL01_CLR1_n_864);
  TL01_CLR1_g41149 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_749, A2 => TL01_CLR1_n_404, B1 => TL01_CLR1_n_678, B2 => TL01_CLR1_n_580, ZN => TL01_CLR1_n_863);
  TL01_CLR1_g41150 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_659, A2 => TL01_CLR1_n_665, B1 => TL01_CLR1_n_461, B2 => TL01_CLR1_n_101, ZN => TL01_CLR1_n_862);
  TL01_CLR1_g41151 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_655, A2 => TL01_CLR1_n_668, B1 => TL01_CLR1_n_459, B2 => TL01_CLR1_n_101, ZN => TL01_CLR1_n_861);
  TL01_CLR1_g41152 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_742, A2 => TL01_CLR1_n_330, B1 => TL01_CLR1_n_622, B2 => TL01_CLR1_n_394, ZN => TL01_CLR1_n_860);
  TL01_CLR1_g41153 : AO22D0BWP7T port map(A1 => TL01_CLR1_n_770, A2 => TL01_CLR1_n_494, B1 => TL01_CLR1_n_491, B2 => TL01_CLR1_n_763, Z => TL01_CLR1_n_859);
  TL01_CLR1_g41154 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_742, A2 => TL01_CLR1_n_412, B1 => TL01_CLR1_n_675, B2 => TL01_CLR1_n_307, ZN => TL01_CLR1_n_858);
  TL01_CLR1_g41155 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_741, A2 => TL01_CLR1_n_368, B1 => TL01_CLR1_n_642, B2 => TL01_CLR1_n_622, ZN => TL01_CLR1_n_857);
  TL01_CLR1_g41156 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_747, A2 => TL01_CLR1_n_405, B1 => TL01_CLR1_n_721, B2 => TL01_CLR1_n_368, ZN => TL01_CLR1_n_856);
  TL01_CLR1_g41157 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_676, A2 => TL01_CLR1_n_486, B1 => TL01_CLR1_n_743, B2 => TL01_CLR1_n_602, ZN => TL01_CLR1_n_855);
  TL01_CLR1_g41158 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_721, A2 => TL01_CLR1_n_745, B1 => TL01_CLR1_n_747, B2 => TL01_CLR1_n_288, ZN => TL01_CLR1_n_854);
  TL01_CLR1_g41159 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_749, A2 => TL01_CLR1_n_323, B1 => TL01_CLR1_n_743, B2 => TL01_CLR1_n_236, ZN => TL01_CLR1_n_853);
  TL01_CLR1_g41160 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_741, A2 => TL01_CLR1_n_288, B1 => TL01_CLR1_n_679, B2 => TL01_CLR1_n_406, ZN => TL01_CLR1_n_852);
  TL01_CLR1_g41161 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_747, A2 => TL01_CLR1_n_398, B1 => TL01_CLR1_n_721, B2 => TL01_CLR1_n_290, ZN => TL01_CLR1_n_851);
  TL01_CLR1_g41162 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_747, A2 => TL01_CLR1_n_306, B1 => TL01_CLR1_n_721, B2 => TL01_CLR1_n_235, ZN => TL01_CLR1_n_850);
  TL01_CLR1_g41163 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_720, A2 => TL01_CLR1_n_732, B => TL01_CLR1_n_812, ZN => TL01_CLR1_n_886);
  TL01_CLR1_g41164 : XNR2D1BWP7T port map(A1 => TL01_CLR1_n_664, A2 => TL01_CLR1_n_458, ZN => TL01_CLR1_n_885);
  TL01_CLR1_g41165 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_663, A2 => TL01_CLR1_n_457, B1 => TL01_CLR1_n_663, B2 => TL01_CLR1_n_457, ZN => TL01_CLR1_n_884);
  TL01_CLR1_g41166 : NR3D0BWP7T port map(A1 => TL01_CLR1_n_746, A2 => TL01_CLR1_n_722, A3 => TL01_CLR1_n_377, ZN => TL01_CLR1_n_883);
  TL01_CLR1_g41167 : INVD0BWP7T port map(I => TL01_CLR1_n_725, ZN => TL01_CLR1_n_849);
  TL01_CLR1_g41168 : INVD1BWP7T port map(I => TL01_CLR1_n_728, ZN => TL01_CLR1_n_848);
  TL01_CLR1_g41169 : INVD0BWP7T port map(I => TL01_CLR1_n_841, ZN => TL01_CLR1_n_842);
  TL01_CLR1_g41170 : INVD0BWP7T port map(I => TL01_CLR1_n_831, ZN => TL01_CLR1_n_832);
  TL01_CLR1_g41171 : INVD0BWP7T port map(I => TL01_CLR1_n_828, ZN => TL01_CLR1_n_829);
  TL01_CLR1_g41172 : INVD0BWP7T port map(I => TL01_CLR1_n_818, ZN => TL01_CLR1_n_817);
  TL01_CLR1_g41173 : INVD0BWP7T port map(I => TL01_CLR1_n_816, ZN => TL01_CLR1_n_815);
  TL01_CLR1_g41174 : INVD0BWP7T port map(I => TL01_CLR1_n_814, ZN => TL01_CLR1_n_813);
  TL01_CLR1_g41175 : INVD1BWP7T port map(I => TL01_CLR1_n_812, ZN => TL01_CLR1_n_811);
  TL01_CLR1_g41176 : NR2D0BWP7T port map(A1 => TL01_CLR1_n_661, A2 => TL01_CLR1_char1_sprite_sprite_0, ZN => TL01_CLR1_n_810);
  TL01_CLR1_g41179 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_717, A2 => TL01_CLR1_n_746, ZN => TL01_CLR1_n_847);
  TL01_CLR1_g41180 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_718, A2 => TL01_CLR1_n_621, ZN => TL01_CLR1_n_846);
  TL01_CLR1_g41181 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_772, A2 => TL01_CLR1_n_456, ZN => TL01_CLR1_n_845);
  TL01_CLR1_g41182 : INR2XD0BWP7T port map(A1 => TL01_CLR1_n_559, B1 => TL01_CLR1_n_749, ZN => TL01_CLR1_n_844);
  TL01_CLR1_g41183 : NR2D0BWP7T port map(A1 => TL01_CLR1_n_741, A2 => TL01_CLR1_n_486, ZN => TL01_CLR1_n_843);
  TL01_CLR1_g41184 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_740, A2 => TL01_CLR1_n_582, ZN => TL01_CLR1_n_841);
  TL01_CLR1_g41185 : INR2D0BWP7T port map(A1 => TL01_CLR1_n_732, B1 => TL01_CLR1_n_718, ZN => TL01_CLR1_n_840);
  TL01_CLR1_g41186 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_742, A2 => TL01_CLR1_n_746, ZN => TL01_CLR1_n_839);
  TL01_CLR1_g41187 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_747, A2 => TL01_CLR1_n_724, ZN => TL01_CLR1_n_838);
  TL01_CLR1_g41188 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_771, A2 => TL01_CLR1_n_158, ZN => TL01_CLR1_n_837);
  TL01_CLR1_g41189 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_717, A2 => TL01_CLR1_n_308, ZN => TL01_CLR1_n_836);
  TL01_CLR1_g41190 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_639, A2 => char1posy(5), ZN => TL01_CLR1_n_835);
  TL01_CLR1_g41191 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_723, A2 => hcountintern(4), ZN => TL01_CLR1_n_834);
  TL01_CLR1_g41192 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_635, A2 => char2posy(5), ZN => TL01_CLR1_n_833);
  TL01_CLR1_g41193 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_720, A2 => TL01_CLR1_n_404, ZN => TL01_CLR1_n_831);
  TL01_CLR1_g41194 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_731, A2 => char2perc(0), ZN => TL01_CLR1_n_830);
  TL01_CLR1_g41195 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_740, A2 => TL01_CLR1_n_283, ZN => TL01_CLR1_n_828);
  TL01_CLR1_g41196 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_662, A2 => TL01_CLR1_char2_sprite_sprite_0, ZN => TL01_CLR1_n_827);
  TL01_CLR1_g41197 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_637, A2 => char1posx(5), ZN => TL01_CLR1_n_826);
  TL01_CLR1_g41198 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_718, A2 => TL01_CLR1_n_237, ZN => TL01_CLR1_n_825);
  TL01_CLR1_g41199 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_641, A2 => char2posx(5), ZN => TL01_CLR1_n_824);
  TL01_CLR1_g41200 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_755, A2 => TL01_CLR1_n_578, ZN => TL01_CLR1_n_823);
  TL01_CLR1_g41201 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_717, A2 => TL01_CLR1_n_675, ZN => TL01_CLR1_n_822);
  TL01_CLR1_g41202 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_744, A2 => TL01_CLR1_n_676, ZN => TL01_CLR1_n_821);
  TL01_CLR1_g41203 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_740, A2 => TL01_CLR1_n_717, ZN => TL01_CLR1_n_820);
  TL01_CLR1_g41204 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_747, A2 => TL01_CLR1_n_721, ZN => TL01_CLR1_n_819);
  TL01_CLR1_g41205 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_751, A2 => TL01_CLR1_n_512, ZN => TL01_CLR1_n_818);
  TL01_CLR1_g41206 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_754, A2 => TL01_CLR1_n_718, ZN => TL01_CLR1_n_816);
  TL01_CLR1_g41207 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_739, A2 => TL01_CLR1_n_600, ZN => TL01_CLR1_n_814);
  TL01_CLR1_g41208 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_754, A2 => TL01_CLR1_n_721, ZN => TL01_CLR1_n_812);
  TL01_CLR1_g41209 : INVD0BWP7T port map(I => TL01_CLR1_n_806, ZN => TL01_CLR1_n_805);
  TL01_CLR1_g41210 : INVD1BWP7T port map(I => TL01_CLR1_n_801, ZN => TL01_CLR1_n_800);
  TL01_CLR1_g41211 : INVD1BWP7T port map(I => TL01_CLR1_n_799, ZN => TL01_CLR1_n_798);
  TL01_CLR1_g41212 : AO211D0BWP7T port map(A1 => TL01_CLR1_n_571, A2 => TL01_CLR1_n_395, B => TL01_CLR1_n_667, C => TL01_CLR1_n_159, Z => TL01_CLR1_n_797);
  TL01_CLR1_g41213 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_206, A2 => TL01_CLR1_n_60, B1 => TL01_CLR1_n_1563, B2 => TL01_CLR1_n_167, C => TL01_CLR1_n_706, ZN => TL01_CLR1_n_796);
  TL01_CLR1_g41214 : AOI31D0BWP7T port map(A1 => TL01_CLR1_n_633, A2 => TL01_CLR1_n_397, A3 => TL01_CLR1_n_341, B => TL01_CLR1_n_697, ZN => TL01_CLR1_n_795);
  TL01_CLR1_g41215 : IAO21D0BWP7T port map(A1 => TL01_CLR1_n_124, A2 => TL01_CLR1_n_145, B => TL01_CLR1_n_771, ZN => TL01_CLR1_n_794);
  TL01_CLR1_g41216 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_687, A2 => TL01_CLR1_n_313, B1 => TL01_CLR1_n_559, B2 => TL01_CLR1_n_193, ZN => TL01_CLR1_n_793);
  TL01_CLR1_g41217 : AN3D0BWP7T port map(A1 => TL01_CLR1_n_692, A2 => TL01_CLR1_n_653, A3 => TL01_CLR1_n_147, Z => TL01_CLR1_n_792);
  TL01_CLR1_g41218 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_583, A2 => vcountintern(5), B => TL01_CLR1_n_666, ZN => TL01_CLR1_n_791);
  TL01_CLR1_g41219 : AOI31D0BWP7T port map(A1 => TL01_CLR1_n_571, A2 => TL01_CLR1_n_628, A3 => TL01_CLR1_n_486, B => TL01_CLR1_n_674, ZN => TL01_CLR1_n_790);
  TL01_CLR1_g41220 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_578, A2 => TL01_CLR1_n_487, B => TL01_CLR1_n_748, ZN => TL01_CLR1_n_789);
  TL01_CLR1_g41221 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_673, A2 => TL01_CLR1_n_321, B1 => TL01_CLR1_n_561, B2 => TL01_CLR1_n_406, ZN => TL01_CLR1_n_788);
  TL01_CLR1_g41222 : ND4D0BWP7T port map(A1 => TL01_CLR1_n_740, A2 => TL01_CLR1_n_309, A3 => TL01_CLR1_n_238, A4 => TL01_CLR1_n_1495, ZN => TL01_CLR1_n_787);
  TL01_CLR1_g41223 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_44, A2 => TL01_CLR1_n_322, B1 => TL01_CLR1_n_561, B2 => TL01_CLR1_n_193, ZN => TL01_CLR1_n_786);
  TL01_CLR1_g41224 : NR4D0BWP7T port map(A1 => TL01_CLR1_n_614, A2 => TL01_CLR1_n_1494, A3 => TL01_CLR1_n_166, A4 => vcountintern(6), ZN => TL01_CLR1_n_785);
  TL01_CLR1_g41225 : NR3D0BWP7T port map(A1 => TL01_CLR1_n_654, A2 => TL01_CLR1_n_625, A3 => TL01_CLR1_n_627, ZN => TL01_CLR1_n_784);
  TL01_CLR1_g41226 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_684, A2 => TL01_CLR1_n_318, B => TL01_CLR1_n_749, ZN => TL01_CLR1_n_783);
  TL01_CLR1_g41227 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_367, A2 => TL01_CLR1_n_308, B => TL01_CLR1_n_717, ZN => TL01_CLR1_n_782);
  TL01_CLR1_g41228 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_498, A2 => TL01_CLR1_n_395, B => TL01_CLR1_n_741, ZN => TL01_CLR1_n_781);
  TL01_CLR1_g41229 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_171, A2 => TL01_CLR1_n_421, B => TL01_CLR1_n_657, C => TL01_CLR1_n_534, ZN => TL01_CLR1_n_780);
  TL01_CLR1_g41230 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_44, A2 => TL01_CLR1_n_495, B1 => TL01_CLR1_n_561, B2 => TL01_CLR1_n_490, ZN => TL01_CLR1_n_779);
  TL01_CLR1_g41231 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_44, A2 => TL01_CLR1_n_403, B1 => TL01_CLR1_n_561, B2 => TL01_CLR1_n_320, ZN => TL01_CLR1_n_778);
  TL01_CLR1_g41232 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_677, A2 => TL01_CLR1_n_285, B1 => TL01_CLR1_n_678, B2 => TL01_CLR1_n_323, ZN => TL01_CLR1_n_777);
  TL01_CLR1_g41233 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_679, A2 => TL01_CLR1_n_314, B1 => TL01_CLR1_n_673, B2 => TL01_CLR1_n_491, ZN => TL01_CLR1_n_776);
  TL01_CLR1_g41234 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_687, A2 => TL01_CLR1_n_314, B1 => TL01_CLR1_n_577, B2 => TL01_CLR1_n_327, ZN => TL01_CLR1_n_775);
  TL01_CLR1_g41235 : AO22D0BWP7T port map(A1 => TL01_CLR1_n_675, A2 => TL01_CLR1_n_408, B1 => TL01_CLR1_n_334, B2 => TL01_CLR1_n_678, Z => TL01_CLR1_n_774);
  TL01_CLR1_g41236 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_685, A2 => TL01_CLR1_n_684, B1 => TL01_CLR1_n_687, B2 => TL01_CLR1_n_198, ZN => TL01_CLR1_n_773);
  TL01_CLR1_g41237 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_569, A2 => char1posx(5), B => TL01_CLR1_n_758, ZN => TL01_CLR1_n_809);
  TL01_CLR1_g41238 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_326, A2 => TL01_CLR1_n_349, B => TL01_CLR1_n_699, ZN => TL01_CLR1_n_808);
  TL01_CLR1_g41239 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_567, A2 => char2posx(5), B => TL01_CLR1_n_760, ZN => TL01_CLR1_n_807);
  TL01_CLR1_g41240 : ND4D0BWP7T port map(A1 => TL01_CLR1_n_691, A2 => TL01_CLR1_n_361, A3 => TL01_CLR1_n_205, A4 => TL01_CLR1_n_158, ZN => TL01_CLR1_n_806);
  TL01_CLR1_g41241 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_568, A2 => char1posy(5), B1 => TL01_CLR1_n_568, B2 => char1posy(5), ZN => TL01_CLR1_n_804);
  TL01_CLR1_g41242 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_570, A2 => char2posy(5), B1 => TL01_CLR1_n_570, B2 => char2posy(5), ZN => TL01_CLR1_n_803);
  TL01_CLR1_g41243 : IOA21D1BWP7T port map(A1 => TL01_CLR1_n_693, A2 => TL01_CLR1_n_504, B => TL01_CLR1_n_724, ZN => TL01_CLR1_n_802);
  TL01_CLR1_g41244 : AOI211XD0BWP7T port map(A1 => TL01_CLR1_n_173, A2 => TL01_CLR1_n_120, B => TL01_CLR1_n_702, C => TL01_CLR1_n_536, ZN => TL01_CLR1_n_801);
  TL01_CLR1_g41245 : NR3D0BWP7T port map(A1 => TL01_CLR1_n_667, A2 => TL01_CLR1_n_209, A3 => TL01_CLR1_n_114, ZN => TL01_CLR1_n_799);
  TL01_CLR1_g41246 : INVD0BWP7T port map(I => TL01_CLR1_n_661, ZN => TL01_CLR1_n_772);
  TL01_CLR1_g41247 : CKND1BWP7T port map(I => TL01_CLR1_n_765, ZN => TL01_CLR1_n_766);
  TL01_CLR1_g41248 : INVD1BWP7T port map(I => TL01_CLR1_n_760, ZN => TL01_CLR1_n_761);
  TL01_CLR1_g41249 : INVD1BWP7T port map(I => TL01_CLR1_n_756, ZN => TL01_CLR1_n_755);
  TL01_CLR1_g41250 : INVD0BWP7T port map(I => TL01_CLR1_n_754, ZN => TL01_CLR1_n_753);
  TL01_CLR1_g41251 : INVD0BWP7T port map(I => TL01_CLR1_n_751, ZN => TL01_CLR1_n_750);
  TL01_CLR1_g41252 : INVD0BWP7T port map(I => TL01_CLR1_n_749, ZN => TL01_CLR1_n_748);
  TL01_CLR1_g41253 : INVD1BWP7T port map(I => TL01_CLR1_n_746, ZN => TL01_CLR1_n_745);
  TL01_CLR1_g41254 : INVD1BWP7T port map(I => TL01_CLR1_n_744, ZN => TL01_CLR1_n_743);
  TL01_CLR1_g41255 : INVD1BWP7T port map(I => TL01_CLR1_n_742, ZN => TL01_CLR1_n_741);
  TL01_CLR1_g41256 : INVD1BWP7T port map(I => TL01_CLR1_n_740, ZN => TL01_CLR1_n_739);
  TL01_CLR1_g41257 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_677, A2 => TL01_CLR1_n_688, ZN => TL01_CLR1_n_738);
  TL01_CLR1_g41258 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_474, A2 => TL01_CLR1_n_1483, B1 => FE_PHN147_TL01_CLR1_n_257, B2 => TL01_CLR1_n_372, C => TL01_CLR1_n_648, ZN => TL01_CLR1_n_737);
  TL01_CLR1_g41259 : ND2D0BWP7T port map(A1 => TL01_CLR1_n_689, A2 => TL01_CLR1_n_623, ZN => TL01_CLR1_n_736);
  TL01_CLR1_g41260 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_649, A2 => TL01_CLR1_n_617, ZN => TL01_CLR1_n_735);
  TL01_CLR1_g41261 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_684, A2 => TL01_CLR1_n_323, Z => TL01_CLR1_n_734);
  TL01_CLR1_g41262 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_480, A2 => TL01_CLR1_char1_sprite_frame_control_state_1, B1 => TL01_CLR1_n_1492, B2 => TL01_CLR1_n_466, C => TL01_CLR1_n_647, ZN => TL01_CLR1_n_733);
  TL01_CLR1_g41263 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_691, A2 => TL01_CLR1_n_166, ZN => TL01_CLR1_n_771);
  TL01_CLR1_g41264 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_624, B1 => TL01_CLR1_n_679, ZN => TL01_CLR1_n_770);
  TL01_CLR1_g41265 : NR3D0BWP7T port map(A1 => TL01_CLR1_n_607, A2 => TL01_CLR1_n_527, A3 => hcountintern(9), ZN => TL01_CLR1_n_769);
  TL01_CLR1_g41266 : ND2D0BWP7T port map(A1 => TL01_CLR1_n_697, A2 => TL01_CLR1_n_399, ZN => TL01_CLR1_n_768);
  TL01_CLR1_g41267 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_677, A2 => TL01_CLR1_n_318, ZN => TL01_CLR1_n_767);
  TL01_CLR1_g41268 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_676, A2 => TL01_CLR1_n_375, ZN => TL01_CLR1_n_765);
  TL01_CLR1_g41269 : NR2D0BWP7T port map(A1 => TL01_CLR1_n_676, A2 => TL01_CLR1_n_487, ZN => TL01_CLR1_n_764);
  TL01_CLR1_g41270 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_686, A2 => TL01_CLR1_n_485, ZN => TL01_CLR1_n_763);
  TL01_CLR1_g41271 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_570, B1 => char2posy(5), ZN => TL01_CLR1_n_762);
  TL01_CLR1_g41272 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_567, A2 => char2posx(5), ZN => TL01_CLR1_n_760);
  TL01_CLR1_g41273 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_568, B1 => char1posy(5), ZN => TL01_CLR1_n_759);
  TL01_CLR1_g41274 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_569, A2 => char1posx(5), ZN => TL01_CLR1_n_758);
  TL01_CLR1_g41275 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_471, A2 => TL01_CLR1_n_300, B1 => TL01_CLR1_n_242, B2 => TL01_CLR1_n_469, C => TL01_CLR1_n_660, ZN => TL01_CLR1_n_757);
  TL01_CLR1_g41276 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_690, A2 => TL01_CLR1_n_492, ZN => TL01_CLR1_n_756);
  TL01_CLR1_g41277 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_693, A2 => TL01_CLR1_n_500, ZN => TL01_CLR1_n_754);
  TL01_CLR1_g41278 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_674, A2 => TL01_CLR1_n_600, ZN => TL01_CLR1_n_752);
  TL01_CLR1_g41279 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_42, A2 => TL01_CLR1_n_410, ZN => TL01_CLR1_n_751);
  TL01_CLR1_g41280 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_561, A2 => TL01_CLR1_n_679, ZN => TL01_CLR1_n_749);
  TL01_CLR1_g41281 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_693, A2 => TL01_CLR1_n_499, ZN => TL01_CLR1_n_747);
  TL01_CLR1_g41282 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_694, A2 => TL01_CLR1_n_200, ZN => TL01_CLR1_n_746);
  TL01_CLR1_g41283 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_688, A2 => vcountintern(0), ZN => TL01_CLR1_n_744);
  TL01_CLR1_g41284 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_689, A2 => vcountintern(0), ZN => TL01_CLR1_n_742);
  TL01_CLR1_g41285 : INR2D1BWP7T port map(A1 => TL01_CLR1_n_693, B1 => TL01_CLR1_n_497, ZN => TL01_CLR1_n_740);
  TL01_CLR1_g41286 : INVD0BWP7T port map(I => TL01_CLR1_n_731, ZN => TL01_CLR1_n_730);
  TL01_CLR1_g41288 : INVD0BWP7T port map(I => TL01_CLR1_n_727, ZN => TL01_CLR1_n_726);
  TL01_CLR1_g41289 : INVD1BWP7T port map(I => TL01_CLR1_n_723, ZN => TL01_CLR1_n_722);
  TL01_CLR1_g41290 : INVD1BWP7T port map(I => TL01_CLR1_n_720, ZN => TL01_CLR1_n_719);
  TL01_CLR1_g41291 : INVD1BWP7T port map(I => TL01_CLR1_n_718, ZN => TL01_CLR1_n_717);
  TL01_CLR1_g41292 : OAI222D0BWP7T port map(A1 => TL01_CLR1_n_556, A2 => TL01_CLR1_n_396, B1 => TL01_CLR1_n_326, B2 => TL01_CLR1_n_397, C1 => TL01_CLR1_n_348, C2 => TL01_CLR1_n_401, ZN => TL01_CLR1_n_716);
  TL01_CLR1_g41293 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_537, A2 => char1perc(1), B1 => TL01_CLR1_n_550, B2 => FE_DBTN13_char1perc_5, C1 => TL01_CLR1_n_555, C2 => char1perc(5), ZN => TL01_CLR1_n_715);
  TL01_CLR1_g41294 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_538, A2 => char1perc(1), B1 => TL01_CLR1_n_441, B2 => TL01_CLR1_n_239, C => TL01_CLR1_n_589, ZN => TL01_CLR1_n_714);
  TL01_CLR1_g41295 : OAI31D0BWP7T port map(A1 => TL01_CLR1_n_248, A2 => TL01_CLR1_n_389, A3 => TL01_CLR1_n_414, B => TL01_CLR1_n_690, ZN => TL01_CLR1_n_713);
  TL01_CLR1_g41296 : AOI211XD0BWP7T port map(A1 => TL01_CLR1_n_399, A2 => TL01_CLR1_n_484, B => TL01_CLR1_n_43, C => TL01_CLR1_n_613, ZN => TL01_CLR1_n_712);
  TL01_CLR1_g41297 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_546, A2 => TL01_CLR1_n_396, B1 => TL01_CLR1_n_644, B2 => TL01_CLR1_n_349, ZN => TL01_CLR1_n_711);
  TL01_CLR1_g41298 : OA222D0BWP7T port map(A1 => TL01_CLR1_n_609, A2 => hcountintern(2), B1 => char1posx(0), B2 => TL01_CLR1_n_66, C1 => char1posx(1), C2 => TL01_CLR1_n_69, Z => TL01_CLR1_n_710);
  TL01_CLR1_g41299 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_505, A2 => TL01_CLR1_n_174, B1 => TL01_CLR1_n_380, B2 => TL01_CLR1_n_419, C => TL01_CLR1_n_645, ZN => TL01_CLR1_n_709);
  TL01_CLR1_g41300 : OAI211D1BWP7T port map(A1 => FE_DBTN12_char1perc_4, A2 => TL01_CLR1_n_521, B => TL01_CLR1_n_360, C => TL01_CLR1_n_354, ZN => TL01_CLR1_n_708);
  TL01_CLR1_g41301 : IAO21D0BWP7T port map(A1 => TL01_CLR1_n_565, A2 => TL01_CLR1_n_197, B => TL01_CLR1_n_686, ZN => TL01_CLR1_n_707);
  TL01_CLR1_g41302 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_531, A2 => TL01_CLR1_n_148, B1 => TL01_CLR1_n_535, B2 => vcountintern(9), C1 => TL01_CLR1_n_271, C2 => TL01_CLR1_n_166, ZN => TL01_CLR1_n_706);
  TL01_CLR1_g41303 : OA222D0BWP7T port map(A1 => TL01_CLR1_n_608, A2 => hcountintern(2), B1 => char2posx(0), B2 => FE_DBTN1_char2posx_1, C1 => char2posx(1), C2 => FE_DBTN0_char2posx_0, Z => TL01_CLR1_n_705);
  TL01_CLR1_g41304 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_590, A2 => TL01_CLR1_n_259, B1 => TL01_CLR1_n_370, B2 => TL01_CLR1_n_1492, ZN => TL01_CLR1_n_704);
  TL01_CLR1_g41305 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_586, A2 => FE_PHN147_TL01_CLR1_n_257, B1 => TL01_CLR1_n_372, B2 => TL01_CLR1_n_1483, ZN => TL01_CLR1_n_703);
  TL01_CLR1_g41306 : OAI221D0BWP7T port map(A1 => TL01_CLR1_n_483, A2 => TL01_CLR1_n_77, B1 => char2perc(7), B2 => TL01_CLR1_n_523, C => TL01_CLR1_n_227, ZN => TL01_CLR1_n_702);
  TL01_CLR1_g41307 : MAOI222D1BWP7T port map(A => TL01_CLR1_n_591, B => TL01_CLR1_n_475, C => TL01_CLR1_n_52, ZN => TL01_CLR1_n_701);
  TL01_CLR1_g41308 : OA21D0BWP7T port map(A1 => TL01_CLR1_n_574, A2 => TL01_CLR1_n_408, B => TL01_CLR1_n_673, Z => TL01_CLR1_n_700);
  TL01_CLR1_g41309 : AO31D1BWP7T port map(A1 => TL01_CLR1_n_573, A2 => TL01_CLR1_n_487, A3 => TL01_CLR1_n_395, B => TL01_CLR1_n_348, Z => TL01_CLR1_n_699);
  TL01_CLR1_g41310 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_543, A2 => TL01_CLR1_n_291, B => TL01_CLR1_n_319, ZN => TL01_CLR1_n_732);
  TL01_CLR1_g41311 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_592, A2 => TL01_CLR1_n_584, A3 => TL01_CLR1_n_594, ZN => TL01_CLR1_n_731);
  TL01_CLR1_g41312 : AOI221D0BWP7T port map(A1 => TL01_CLR1_n_550, A2 => TL01_CLR1_n_175, B1 => TL01_CLR1_n_472, B2 => TL01_CLR1_n_342, C => TL01_CLR1_n_598, ZN => TL01_CLR1_n_729);
  TL01_CLR1_g41313 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_604, A2 => hcountintern(3), B1 => TL01_CLR1_n_604, B2 => hcountintern(3), ZN => TL01_CLR1_n_728);
  TL01_CLR1_g41314 : OAI31D0BWP7T port map(A1 => TL01_CLR1_n_127, A2 => TL01_CLR1_n_102, A3 => TL01_CLR1_n_140, B => TL01_CLR1_n_646, ZN => TL01_CLR1_n_727);
  TL01_CLR1_g41315 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_1561, A2 => hcountintern(3), B1 => TL01_CLR1_n_1561, B2 => hcountintern(3), ZN => TL01_CLR1_n_725);
  TL01_CLR1_g41316 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_633, A2 => TL01_CLR1_n_504, A3 => TL01_CLR1_n_397, ZN => TL01_CLR1_n_724);
  TL01_CLR1_g41317 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_543, A2 => TL01_CLR1_n_200, A3 => TL01_CLR1_n_291, ZN => TL01_CLR1_n_723);
  TL01_CLR1_g41318 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_633, A2 => TL01_CLR1_n_499, A3 => TL01_CLR1_n_52, ZN => TL01_CLR1_n_721);
  TL01_CLR1_g41319 : NR3D0BWP7T port map(A1 => TL01_CLR1_n_549, A2 => TL01_CLR1_n_289, A3 => TL01_CLR1_n_200, ZN => TL01_CLR1_n_720);
  TL01_CLR1_g41320 : ND3D1BWP7T port map(A1 => TL01_CLR1_n_633, A2 => TL01_CLR1_n_500, A3 => TL01_CLR1_n_52, ZN => TL01_CLR1_n_718);
  TL01_CLR1_g41321 : INVD1BWP7T port map(I => TL01_CLR1_n_689, ZN => TL01_CLR1_n_688);
  TL01_CLR1_g41322 : INVD0BWP7T port map(I => TL01_CLR1_n_686, ZN => TL01_CLR1_n_685);
  TL01_CLR1_g41323 : INVD1BWP7T port map(I => TL01_CLR1_n_683, ZN => TL01_CLR1_n_682);
  TL01_CLR1_g41324 : INVD1BWP7T port map(I => TL01_CLR1_n_681, ZN => TL01_CLR1_n_680);
  TL01_CLR1_g41325 : INVD0BWP7T port map(I => TL01_CLR1_n_679, ZN => TL01_CLR1_n_678);
  TL01_CLR1_g41326 : INVD1BWP7T port map(I => TL01_CLR1_n_677, ZN => TL01_CLR1_n_676);
  TL01_CLR1_g41327 : INVD1BWP7T port map(I => TL01_CLR1_n_675, ZN => TL01_CLR1_n_674);
  TL01_CLR1_g41328 : INVD1BWP7T port map(I => TL01_CLR1_n_44, ZN => TL01_CLR1_n_673);
  TL01_CLR1_g41329 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_259, A2 => TL01_CLR1_n_452, B => TL01_CLR1_n_588, C => TL01_CLR1_n_479, ZN => TL01_CLR1_n_672);
  TL01_CLR1_g41330 : OAI211D1BWP7T port map(A1 => FE_PHN147_TL01_CLR1_n_257, A2 => TL01_CLR1_n_449, B => TL01_CLR1_n_587, C => TL01_CLR1_n_453, ZN => TL01_CLR1_n_671);
  TL01_CLR1_g41331 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_496, B1 => TL01_CLR1_n_1493, ZN => TL01_CLR1_n_670);
  TL01_CLR1_g41333 : NR2D0BWP7T port map(A1 => TL01_CLR1_n_621, A2 => TL01_CLR1_n_237, ZN => TL01_CLR1_n_698);
  TL01_CLR1_g41334 : NR3D0BWP7T port map(A1 => TL01_CLR1_n_473, A2 => TL01_CLR1_n_159, A3 => vcountintern(0), ZN => TL01_CLR1_n_697);
  TL01_CLR1_g41335 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_424, A2 => char2posx(0), B => TL01_CLR1_n_509, ZN => TL01_CLR1_n_696);
  TL01_CLR1_g41336 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_418, A2 => char2posy(4), B => TL01_CLR1_n_634, ZN => TL01_CLR1_n_695);
  TL01_CLR1_g41337 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_291, B1 => TL01_CLR1_n_543, ZN => TL01_CLR1_n_694);
  TL01_CLR1_g41338 : NR3D0BWP7T port map(A1 => TL01_CLR1_n_560, A2 => TL01_CLR1_n_396, A3 => vcountintern(0), ZN => TL01_CLR1_n_693);
  TL01_CLR1_g41340 : IOA21D1BWP7T port map(A1 => TL01_CLR1_n_551, A2 => TL01_CLR1_n_68, B => TL01_CLR1_n_147, ZN => TL01_CLR1_n_692);
  TL01_CLR1_g41341 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_615, A2 => TL01_CLR1_n_148, ZN => TL01_CLR1_n_691);
  TL01_CLR1_g41342 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_77, A2 => TL01_CLR1_n_161, B => TL01_CLR1_n_526, C => TL01_CLR1_n_296, ZN => TL01_CLR1_n_690);
  TL01_CLR1_g41343 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_625, A2 => TL01_CLR1_n_349, ZN => TL01_CLR1_n_689);
  TL01_CLR1_g41344 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_620, A2 => TL01_CLR1_n_564, ZN => TL01_CLR1_n_687);
  TL01_CLR1_g41345 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_620, A2 => TL01_CLR1_n_557, ZN => TL01_CLR1_n_686);
  TL01_CLR1_g41346 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_507, A2 => TL01_CLR1_n_314, ZN => TL01_CLR1_n_684);
  TL01_CLR1_g41347 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_627, A2 => vcountintern(1), ZN => TL01_CLR1_n_683);
  TL01_CLR1_g41348 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_600, A2 => TL01_CLR1_n_558, ZN => TL01_CLR1_n_681);
  TL01_CLR1_g41349 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_348, B1 => TL01_CLR1_n_627, ZN => TL01_CLR1_n_679);
  TL01_CLR1_g41350 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_643, A2 => vcountintern(0), ZN => TL01_CLR1_n_677);
  TL01_CLR1_g41351 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_623, A2 => vcountintern(0), ZN => TL01_CLR1_n_675);
  TL01_CLR1_g41353 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_544, A2 => TL01_CLR1_n_174, B1 => TL01_CLR1_n_427, B2 => TL01_CLR1_n_343, C1 => TL01_CLR1_n_419, C2 => TL01_CLR1_n_251, ZN => TL01_CLR1_n_660);
  TL01_CLR1_g41354 : AO21D0BWP7T port map(A1 => TL01_CLR1_n_461, A2 => hcountintern(4), B => hcountintern(5), Z => TL01_CLR1_n_659);
  TL01_CLR1_g41355 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_484, A2 => TL01_CLR1_n_287, B1 => TL01_CLR1_n_559, B2 => TL01_CLR1_n_306, ZN => TL01_CLR1_n_658);
  TL01_CLR1_g41356 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_548, A2 => TL01_CLR1_n_298, B => TL01_CLR1_n_155, ZN => TL01_CLR1_n_657);
  TL01_CLR1_g41357 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_559, A2 => TL01_CLR1_n_398, B1 => TL01_CLR1_n_405, B2 => TL01_CLR1_n_485, ZN => TL01_CLR1_n_656);
  TL01_CLR1_g41358 : AO21D0BWP7T port map(A1 => TL01_CLR1_n_459, A2 => hcountintern(4), B => hcountintern(5), Z => TL01_CLR1_n_655);
  TL01_CLR1_g41359 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_574, A2 => TL01_CLR1_n_488, B1 => TL01_CLR1_n_209, B2 => TL01_CLR1_n_55, ZN => TL01_CLR1_n_654);
  TL01_CLR1_g41360 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_416, A2 => TL01_CLR1_n_86, B => TL01_CLR1_n_1494, ZN => TL01_CLR1_n_653);
  TL01_CLR1_g41361 : AO211D0BWP7T port map(A1 => TL01_CLR1_n_482, A2 => TL01_CLR1_n_112, B => TL01_CLR1_n_505, C => TL01_CLR1_n_425, Z => TL01_CLR1_n_652);
  TL01_CLR1_g41362 : AO21D0BWP7T port map(A1 => TL01_CLR1_n_399, A2 => TL01_CLR1_n_327, B => TL01_CLR1_n_595, Z => TL01_CLR1_n_651);
  TL01_CLR1_g41363 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_562, A2 => TL01_CLR1_n_404, B => TL01_CLR1_n_624, ZN => TL01_CLR1_n_650);
  TL01_CLR1_g41364 : AOI32D1BWP7T port map(A1 => TL01_CLR1_n_434, A2 => TL01_CLR1_n_447, A3 => char1posy(0), B1 => TL01_CLR1_n_481, B2 => vcountintern(2), ZN => TL01_CLR1_n_649);
  TL01_CLR1_g41365 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_540, A2 => TL01_CLR1_n_1480, B1 => TL01_CLR1_n_362, B2 => TL01_CLR1_n_329, ZN => TL01_CLR1_n_648);
  TL01_CLR1_g41366 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_530, A2 => TL01_CLR1_n_1489, B1 => TL01_CLR1_n_370, B2 => TL01_CLR1_n_259, ZN => TL01_CLR1_n_647);
  TL01_CLR1_g41367 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_525, A2 => char2perc(4), B1 => TL01_CLR1_n_296, B2 => TL01_CLR1_n_61, ZN => TL01_CLR1_n_646);
  TL01_CLR1_g41368 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_533, A2 => char2perc(1), B1 => TL01_CLR1_n_437, B2 => TL01_CLR1_n_242, ZN => TL01_CLR1_n_645);
  TL01_CLR1_g41369 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_423, A2 => char1posx(0), B => TL01_CLR1_n_462, ZN => TL01_CLR1_n_669);
  TL01_CLR1_g41370 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_423, A2 => char1posx(4), B => TL01_CLR1_n_636, ZN => TL01_CLR1_n_668);
  TL01_CLR1_g41371 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_416, A2 => vcountintern(4), B1 => TL01_CLR1_n_416, B2 => vcountintern(4), ZN => TL01_CLR1_n_667);
  TL01_CLR1_g41372 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_420, A2 => char1posy(4), B => TL01_CLR1_n_638, ZN => TL01_CLR1_n_666);
  TL01_CLR1_g41373 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_424, A2 => char2posx(4), B => TL01_CLR1_n_640, ZN => TL01_CLR1_n_665);
  TL01_CLR1_g41374 : MAOI222D1BWP7T port map(A => TL01_CLR1_n_542, B => TL01_CLR1_n_1562, C => vcountintern(3), ZN => TL01_CLR1_n_664);
  TL01_CLR1_g41375 : MAOI222D1BWP7T port map(A => TL01_CLR1_n_503, B => TL01_CLR1_n_204, C => vcountintern(3), ZN => TL01_CLR1_n_663);
  TL01_CLR1_g41376 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_503, A2 => TL01_CLR1_n_467, B1 => TL01_CLR1_n_503, B2 => TL01_CLR1_n_467, ZN => TL01_CLR1_n_662);
  TL01_CLR1_g41377 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_542, A2 => TL01_CLR1_n_465, B1 => TL01_CLR1_n_542, B2 => TL01_CLR1_n_465, ZN => TL01_CLR1_n_661);
  TL01_CLR1_g41379 : INVD0BWP7T port map(I => TL01_CLR1_n_640, ZN => TL01_CLR1_n_641);
  TL01_CLR1_g41380 : CKND1BWP7T port map(I => TL01_CLR1_n_638, ZN => TL01_CLR1_n_639);
  TL01_CLR1_g41381 : INVD1BWP7T port map(I => TL01_CLR1_n_636, ZN => TL01_CLR1_n_637);
  TL01_CLR1_g41382 : INVD0BWP7T port map(I => TL01_CLR1_n_634, ZN => TL01_CLR1_n_635);
  TL01_CLR1_g41383 : INVD1BWP7T port map(I => TL01_CLR1_n_632, ZN => TL01_CLR1_n_631);
  TL01_CLR1_g41384 : INVD1BWP7T port map(I => TL01_CLR1_n_628, ZN => TL01_CLR1_n_629);
  TL01_CLR1_g41385 : INVD0BWP7T port map(I => TL01_CLR1_n_626, ZN => TL01_CLR1_n_625);
  TL01_CLR1_g41386 : INVD1BWP7T port map(I => TL01_CLR1_n_623, ZN => TL01_CLR1_n_622);
  TL01_CLR1_g41387 : INVD1BWP7T port map(I => TL01_CLR1_n_621, ZN => TL01_CLR1_n_620);
  TL01_CLR1_g41388 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_562, B1 => TL01_CLR1_n_375, ZN => TL01_CLR1_n_619);
  TL01_CLR1_g41389 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_396, A2 => TL01_CLR1_n_114, B => TL01_CLR1_n_546, ZN => TL01_CLR1_n_618);
  TL01_CLR1_g41390 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_386, A2 => vcountintern(4), B1 => TL01_CLR1_n_446, B2 => vcountintern(3), ZN => TL01_CLR1_n_617);
  TL01_CLR1_g41391 : OA21D0BWP7T port map(A1 => TL01_CLR1_n_462, A2 => FE_DBTN3_char1posx_4, B => TL01_CLR1_n_569, Z => TL01_CLR1_n_616);
  TL01_CLR1_g41392 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_86, A2 => TL01_CLR1_n_333, B => TL01_CLR1_n_436, C => TL01_CLR1_n_169, ZN => TL01_CLR1_n_615);
  TL01_CLR1_g41393 : OAI211D1BWP7T port map(A1 => hcountintern(7), A2 => TL01_CLR1_n_357, B => TL01_CLR1_n_206, C => TL01_CLR1_n_282, ZN => TL01_CLR1_n_614);
  TL01_CLR1_g41394 : NR2D0BWP7T port map(A1 => TL01_CLR1_n_559, A2 => TL01_CLR1_n_413, ZN => TL01_CLR1_n_613);
  TL01_CLR1_g41395 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_562, A2 => TL01_CLR1_n_307, ZN => TL01_CLR1_n_612);
  TL01_CLR1_g41396 : INR2XD0BWP7T port map(A1 => TL01_CLR1_n_457, B1 => TL01_CLR1_n_1494, ZN => TL01_CLR1_n_611);
  TL01_CLR1_g41397 : CKAN2D1BWP7T port map(A1 => TL01_CLR1_n_573, A2 => TL01_CLR1_n_401, Z => TL01_CLR1_n_644);
  TL01_CLR1_g41398 : OA21D0BWP7T port map(A1 => TL01_CLR1_n_509, A2 => TL01_CLR1_n_75, B => TL01_CLR1_n_567, Z => TL01_CLR1_n_610);
  TL01_CLR1_g41399 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_497, B1 => TL01_CLR1_n_560, ZN => TL01_CLR1_n_643);
  TL01_CLR1_g41400 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_565, A2 => TL01_CLR1_n_286, Z => TL01_CLR1_n_642);
  TL01_CLR1_g41401 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_424, A2 => char2posx(4), ZN => TL01_CLR1_n_640);
  TL01_CLR1_g41402 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_420, A2 => char1posy(4), ZN => TL01_CLR1_n_638);
  TL01_CLR1_g41403 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_423, A2 => char1posx(4), ZN => TL01_CLR1_n_636);
  TL01_CLR1_g41404 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_418, A2 => char2posy(4), ZN => TL01_CLR1_n_634);
  TL01_CLR1_g41405 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_560, A2 => TL01_CLR1_n_55, ZN => TL01_CLR1_n_633);
  TL01_CLR1_g41406 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_77, A2 => TL01_CLR1_n_390, B => TL01_CLR1_n_438, C => TL01_CLR1_n_227, ZN => TL01_CLR1_n_632);
  TL01_CLR1_g41407 : AOI211D1BWP7T port map(A1 => TL01_CLR1_n_240, A2 => TL01_CLR1_n_178, B => TL01_CLR1_n_541, C => TL01_CLR1_n_358, ZN => TL01_CLR1_n_630);
  TL01_CLR1_g41408 : IND3D1BWP7T port map(A1 => TL01_CLR1_n_289, B1 => TL01_CLR1_n_200, B2 => TL01_CLR1_n_460, ZN => TL01_CLR1_n_628);
  TL01_CLR1_g41409 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_473, A2 => TL01_CLR1_n_209, ZN => TL01_CLR1_n_627);
  TL01_CLR1_g41410 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_560, A2 => TL01_CLR1_n_433, ZN => TL01_CLR1_n_626);
  TL01_CLR1_g41411 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_559, A2 => TL01_CLR1_n_485, ZN => TL01_CLR1_n_624);
  TL01_CLR1_g41412 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_560, A2 => TL01_CLR1_n_499, ZN => TL01_CLR1_n_623);
  TL01_CLR1_g41413 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_500, A2 => vcountintern(3), A3 => vcountintern(0), ZN => TL01_CLR1_n_621);
  TL01_CLR1_g41414 : MAOI222D1BWP7T port map(A => TL01_CLR1_n_515, B => TL01_CLR1_n_350, C => hcountintern(3), ZN => TL01_CLR1_n_599);
  TL01_CLR1_g41415 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_443, A2 => TL01_CLR1_n_171, B1 => TL01_CLR1_n_470, B2 => TL01_CLR1_n_240, ZN => TL01_CLR1_n_598);
  TL01_CLR1_g41416 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_463, A2 => TL01_CLR1_n_150, B => TL01_CLR1_n_146, ZN => TL01_CLR1_n_597);
  TL01_CLR1_g41417 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_464, A2 => TL01_CLR1_n_150, B => TL01_CLR1_n_146, ZN => TL01_CLR1_n_596);
  TL01_CLR1_g41418 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_493, A2 => TL01_CLR1_n_413, B => TL01_CLR1_n_563, ZN => TL01_CLR1_n_595);
  TL01_CLR1_g41419 : OA22D0BWP7T port map(A1 => TL01_CLR1_n_471, A2 => TL01_CLR1_n_242, B1 => TL01_CLR1_n_102, B2 => TL01_CLR1_n_297, Z => TL01_CLR1_n_594);
  TL01_CLR1_g41420 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_405, A2 => TL01_CLR1_n_284, B => TL01_CLR1_n_558, ZN => TL01_CLR1_n_593);
  TL01_CLR1_g41421 : AOI32D1BWP7T port map(A1 => TL01_CLR1_n_380, A2 => TL01_CLR1_n_192, A3 => TL01_CLR1_n_174, B1 => TL01_CLR1_n_468, B2 => TL01_CLR1_n_251, ZN => TL01_CLR1_n_592);
  TL01_CLR1_g41422 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_440, A2 => char2posy(0), B1 => TL01_CLR1_n_144, B2 => vcountintern(2), ZN => TL01_CLR1_n_591);
  TL01_CLR1_g41423 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_370, A2 => TL01_CLR1_n_278, B1 => TL01_CLR1_n_466, B2 => inputsp1(3), ZN => TL01_CLR1_n_590);
  TL01_CLR1_g41424 : AOI32D1BWP7T port map(A1 => TL01_CLR1_n_382, A2 => TL01_CLR1_n_170, A3 => TL01_CLR1_n_155, B1 => TL01_CLR1_n_506, B2 => TL01_CLR1_n_175, ZN => TL01_CLR1_n_589);
  TL01_CLR1_g41425 : OA32D1BWP7T port map(A1 => TL01_CLR1_n_1490, A2 => TL01_CLR1_n_338, A3 => TL01_CLR1_n_1489, B1 => TL01_CLR1_n_1492, B2 => TL01_CLR1_n_1484, Z => TL01_CLR1_n_588);
  TL01_CLR1_g41426 : OA32D1BWP7T port map(A1 => TL01_CLR1_n_1481, A2 => TL01_CLR1_n_339, A3 => TL01_CLR1_n_1480, B1 => TL01_CLR1_n_1483, B2 => TL01_CLR1_n_1475, Z => TL01_CLR1_n_587);
  TL01_CLR1_g41427 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_372, A2 => TL01_CLR1_n_279, B1 => TL01_CLR1_n_474, B2 => inputsp2(3), ZN => TL01_CLR1_n_586);
  TL01_CLR1_g41428 : MAOI222D1BWP7T port map(A => TL01_CLR1_n_517, B => TL01_CLR1_n_211, C => hcountintern(3), ZN => TL01_CLR1_n_585);
  TL01_CLR1_g41429 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_505, A2 => TL01_CLR1_n_343, B1 => TL01_CLR1_n_381, B2 => TL01_CLR1_n_419, ZN => TL01_CLR1_n_584);
  TL01_CLR1_g41430 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_463, A2 => TL01_CLR1_n_54, B1 => TL01_CLR1_n_85, B2 => TL01_CLR1_n_69, ZN => TL01_CLR1_n_609);
  TL01_CLR1_g41431 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_464, A2 => TL01_CLR1_n_54, B1 => TL01_CLR1_n_85, B2 => FE_DBTN0_char2posx_0, ZN => TL01_CLR1_n_608);
  TL01_CLR1_g41432 : OR4XD1BWP7T port map(A1 => TL01_CLR1_n_106, A2 => TL01_CLR1_n_1494, A3 => TL01_CLR1_n_148, A4 => TL01_CLR1_n_429, Z => TL01_CLR1_n_607);
  TL01_CLR1_g41433 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_335, A2 => char2posy(4), B1 => TL01_CLR1_n_335, B2 => char2posy(4), ZN => TL01_CLR1_n_606);
  TL01_CLR1_g41435 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_515, A2 => TL01_CLR1_n_212, B1 => TL01_CLR1_n_515, B2 => TL01_CLR1_n_212, ZN => TL01_CLR1_n_604);
  TL01_CLR1_g41436 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_336, A2 => char1posy(4), B1 => TL01_CLR1_n_336, B2 => char1posy(4), ZN => TL01_CLR1_n_603);
  TL01_CLR1_g41437 : AN3D1BWP7T port map(A1 => TL01_CLR1_n_460, A2 => TL01_CLR1_n_289, A3 => TL01_CLR1_n_199, Z => TL01_CLR1_n_602);
  TL01_CLR1_g41438 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_442, A2 => char1perc(4), B => TL01_CLR1_n_532, ZN => TL01_CLR1_n_601);
  TL01_CLR1_g41439 : IND3D1BWP7T port map(A1 => TL01_CLR1_n_209, B1 => TL01_CLR1_n_116, B2 => TL01_CLR1_n_560, ZN => TL01_CLR1_n_600);
  TL01_CLR1_g41440 : CKND1BWP7T port map(I => TL01_CLR1_n_458, ZN => TL01_CLR1_n_583);
  TL01_CLR1_g41441 : INVD0BWP7T port map(I => TL01_CLR1_n_564, ZN => TL01_CLR1_n_563);
  TL01_CLR1_g41442 : INVD1BWP7T port map(I => TL01_CLR1_n_558, ZN => TL01_CLR1_n_557);
  TL01_CLR1_g41443 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_486, A2 => TL01_CLR1_n_349, Z => TL01_CLR1_n_556);
  TL01_CLR1_g41444 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_472, B1 => TL01_CLR1_n_421, ZN => TL01_CLR1_n_555);
  TL01_CLR1_g41445 : ND2D0BWP7T port map(A1 => TL01_CLR1_n_493, A2 => TL01_CLR1_n_288, ZN => TL01_CLR1_n_554);
  TL01_CLR1_g41446 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_463, A2 => TL01_CLR1_n_54, ZN => TL01_CLR1_n_553);
  TL01_CLR1_g41447 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_464, A2 => TL01_CLR1_n_54, ZN => TL01_CLR1_n_552);
  TL01_CLR1_g41448 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_392, A2 => vcountintern(6), B => vcountintern(7), ZN => TL01_CLR1_n_551);
  TL01_CLR1_g41449 : AN2D1BWP7T port map(A1 => TL01_CLR1_n_489, A2 => TL01_CLR1_n_233, Z => TL01_CLR1_n_582);
  TL01_CLR1_g41450 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_497, B1 => TL01_CLR1_n_126, ZN => TL01_CLR1_n_581);
  TL01_CLR1_g41451 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_493, A2 => TL01_CLR1_n_320, ZN => TL01_CLR1_n_580);
  TL01_CLR1_g41452 : AN2D1BWP7T port map(A1 => TL01_CLR1_n_489, A2 => TL01_CLR1_n_320, Z => TL01_CLR1_n_579);
  TL01_CLR1_g41453 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_501, A2 => TL01_CLR1_n_408, ZN => TL01_CLR1_n_578);
  TL01_CLR1_g41454 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_512, A2 => TL01_CLR1_n_310, Z => TL01_CLR1_n_577);
  TL01_CLR1_g41455 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_50, A2 => TL01_CLR1_char1_sprite_sprite_1, ZN => TL01_CLR1_n_576);
  TL01_CLR1_g41456 : ND2D1BWP7T port map(A1 => TL01_CLR1_char1_sprite_sprite_0, A2 => TL01_CLR1_char1_sprite_sprite_1, ZN => TL01_CLR1_n_575);
  TL01_CLR1_g41457 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_498, A2 => TL01_CLR1_n_486, ZN => TL01_CLR1_n_574);
  TL01_CLR1_g41458 : CKAN2D1BWP7T port map(A1 => TL01_CLR1_n_486, A2 => TL01_CLR1_n_326, Z => TL01_CLR1_n_573);
  TL01_CLR1_g41459 : CKAN2D1BWP7T port map(A1 => TL01_CLR1_n_513, A2 => TL01_CLR1_n_1495, Z => TL01_CLR1_n_572);
  TL01_CLR1_g41460 : CKAN2D1BWP7T port map(A1 => TL01_CLR1_n_498, A2 => TL01_CLR1_n_401, Z => TL01_CLR1_n_571);
  TL01_CLR1_g41461 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_335, B1 => char2posy(4), ZN => TL01_CLR1_n_570);
  TL01_CLR1_g41462 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_462, A2 => FE_DBTN3_char1posx_4, ZN => TL01_CLR1_n_569);
  TL01_CLR1_g41463 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_336, B1 => char1posy(4), ZN => TL01_CLR1_n_568);
  TL01_CLR1_g41464 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_509, A2 => TL01_CLR1_n_75, ZN => TL01_CLR1_n_567);
  TL01_CLR1_g41465 : INR2D1BWP7T port map(A1 => TL01_CLR1_char2_sprite_sprite_0, B1 => TL01_CLR1_char2_sprite_sprite_1, ZN => TL01_CLR1_n_566);
  TL01_CLR1_g41466 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_511, A2 => TL01_CLR1_n_311, ZN => TL01_CLR1_n_565);
  TL01_CLR1_g41467 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_497, A2 => TL01_CLR1_n_397, ZN => TL01_CLR1_n_564);
  TL01_CLR1_g41468 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_502, A2 => TL01_CLR1_n_313, ZN => TL01_CLR1_n_562);
  TL01_CLR1_g41469 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_504, A2 => TL01_CLR1_n_126, ZN => TL01_CLR1_n_561);
  TL01_CLR1_g41470 : AO211D0BWP7T port map(A1 => TL01_CLR1_n_52, A2 => TL01_CLR1_n_83, B => TL01_CLR1_n_366, C => TL01_CLR1_n_333, Z => TL01_CLR1_n_560);
  TL01_CLR1_g41471 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_499, A2 => TL01_CLR1_n_126, ZN => TL01_CLR1_n_559);
  TL01_CLR1_g41472 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_500, A2 => TL01_CLR1_n_126, ZN => TL01_CLR1_n_558);
  TL01_CLR1_g41473 : OAI31D0BWP7T port map(A1 => TL01_CLR1_n_56, A2 => FE_DBTN12_char1perc_4, A3 => TL01_CLR1_n_216, B => TL01_CLR1_n_450, ZN => TL01_CLR1_n_541);
  TL01_CLR1_g41474 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_371, A2 => TL01_CLR1_n_1483, B => TL01_CLR1_n_268, ZN => TL01_CLR1_n_540);
  TL01_CLR1_g41475 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_397, A2 => vcountintern(1), B => TL01_CLR1_n_432, ZN => TL01_CLR1_n_539);
  TL01_CLR1_g41476 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_383, A2 => TL01_CLR1_n_228, B1 => TL01_CLR1_n_252, B2 => FE_DBTN12_char1perc_4, ZN => TL01_CLR1_n_538);
  TL01_CLR1_g41477 : AO211D0BWP7T port map(A1 => TL01_CLR1_n_274, A2 => TL01_CLR1_n_110, B => TL01_CLR1_n_506, C => TL01_CLR1_n_299, Z => TL01_CLR1_n_537);
  TL01_CLR1_g41478 : AN3D0BWP7T port map(A1 => TL01_CLR1_n_422, A2 => FE_DBTN9_char2perc_5, A3 => char2perc(4), Z => TL01_CLR1_n_536);
  TL01_CLR1_g41479 : IND4D0BWP7T port map(A1 => vcountintern(8), B1 => TL01_CLR1_n_107, B2 => TL01_CLR1_n_176, B3 => TL01_CLR1_n_295, ZN => TL01_CLR1_n_535);
  TL01_CLR1_g41480 : IND3D1BWP7T port map(A1 => TL01_CLR1_n_191, B1 => TL01_CLR1_n_175, B2 => TL01_CLR1_n_382, ZN => TL01_CLR1_n_534);
  TL01_CLR1_g41481 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_381, A2 => TL01_CLR1_n_391, B1 => TL01_CLR1_n_422, B2 => FE_DBTN8_char2perc_4, ZN => TL01_CLR1_n_533);
  TL01_CLR1_g41482 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_276, A2 => char1perc(4), B1 => TL01_CLR1_n_428, B2 => TL01_CLR1_n_87, ZN => TL01_CLR1_n_532);
  TL01_CLR1_g41483 : AOI211D0BWP7T port map(A1 => TL01_CLR1_n_294, A2 => vcountintern(5), B => TL01_CLR1_n_160, C => TL01_CLR1_n_106, ZN => TL01_CLR1_n_531);
  TL01_CLR1_g41484 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_369, A2 => TL01_CLR1_n_1492, B => TL01_CLR1_n_261, ZN => TL01_CLR1_n_530);
  TL01_CLR1_g41485 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_241, A2 => char2perc(5), B1 => TL01_CLR1_n_161, B2 => TL01_CLR1_n_134, C1 => TL01_CLR1_n_251, C2 => char2perc(1), ZN => TL01_CLR1_n_529);
  TL01_CLR1_g41486 : AOI32D1BWP7T port map(A1 => TL01_CLR1_n_280, A2 => hcountintern(5), A3 => hcountintern(9), B1 => TL01_CLR1_n_205, B2 => TL01_CLR1_n_84, ZN => TL01_CLR1_n_528);
  TL01_CLR1_g41487 : OAI32D1BWP7T port map(A1 => hcountintern(6), A2 => TL01_CLR1_n_82, A3 => TL01_CLR1_n_101, B1 => TL01_CLR1_n_188, B2 => TL01_CLR1_n_356, ZN => TL01_CLR1_n_527);
  TL01_CLR1_g41488 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_275, A2 => char2perc(5), B1 => TL01_CLR1_n_353, B2 => TL01_CLR1_n_61, ZN => TL01_CLR1_n_526);
  TL01_CLR1_g41489 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_121, A2 => char2perc(5), B1 => TL01_CLR1_n_352, B2 => TL01_CLR1_n_120, ZN => TL01_CLR1_n_525);
  TL01_CLR1_g41490 : AOI222D0BWP7T port map(A1 => TL01_CLR1_n_343, A2 => char2perc(7), B1 => TL01_CLR1_n_192, B2 => FE_DBTN5_char2perc_1, C1 => TL01_CLR1_n_174, C2 => TL01_CLR1_n_77, ZN => TL01_CLR1_n_524);
  TL01_CLR1_g41491 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_221, A2 => char2perc(2), B1 => TL01_CLR1_n_390, B2 => FE_DBTN7_char2perc_3, ZN => TL01_CLR1_n_523);
  TL01_CLR1_g41492 : OAI222D0BWP7T port map(A1 => TL01_CLR1_n_196, A2 => char2perc(7), B1 => TL01_CLR1_n_77, B2 => TL01_CLR1_n_172, C1 => FE_DBTN5_char2perc_1, C2 => TL01_CLR1_n_347, ZN => TL01_CLR1_n_522);
  TL01_CLR1_g41493 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_365, A2 => TL01_CLR1_n_56, B1 => TL01_CLR1_n_252, B2 => FE_DBTN13_char1perc_5, ZN => TL01_CLR1_n_521);
  TL01_CLR1_g41494 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_298, A2 => TL01_CLR1_n_156, B1 => TL01_CLR1_n_421, B2 => char1perc(1), ZN => TL01_CLR1_n_520);
  TL01_CLR1_g41495 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_292, A2 => TL01_CLR1_n_152, B => TL01_CLR1_n_444, ZN => TL01_CLR1_n_550);
  TL01_CLR1_g41496 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_258, A2 => hcountintern(3), B => TL01_CLR1_n_507, ZN => TL01_CLR1_n_549);
  TL01_CLR1_g41497 : AO22D0BWP7T port map(A1 => TL01_CLR1_n_383, A2 => TL01_CLR1_n_170, B1 => TL01_CLR1_n_342, B2 => TL01_CLR1_n_240, Z => TL01_CLR1_n_548);
  TL01_CLR1_g41498 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_401, A2 => TL01_CLR1_n_395, A3 => TL01_CLR1_n_238, ZN => TL01_CLR1_n_547);
  TL01_CLR1_g41499 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_414, A2 => TL01_CLR1_n_51, B1 => TL01_CLR1_n_324, B2 => TL01_hcount_int(0), ZN => TL01_CLR1_n_546);
  TL01_CLR1_g41500 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_394, A2 => TL01_CLR1_n_190, A3 => TL01_CLR1_n_55, ZN => TL01_CLR1_n_545);
  TL01_CLR1_g41501 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_293, A2 => TL01_CLR1_n_99, B => TL01_CLR1_n_476, ZN => TL01_CLR1_n_544);
  TL01_CLR1_g41502 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_256, A2 => hcountintern(3), B1 => TL01_CLR1_n_256, B2 => hcountintern(3), ZN => TL01_CLR1_n_543);
  TL01_CLR1_g41503 : OAI211D1BWP7T port map(A1 => char1posy(0), A2 => TL01_CLR1_n_183, B => TL01_CLR1_n_431, C => TL01_CLR1_n_159, ZN => TL01_CLR1_n_542);
  TL01_CLR1_g41504 : INVD0BWP7T port map(I => TL01_CLR1_n_519, ZN => TL01_CLR1_n_518);
  TL01_CLR1_g41505 : CKND1BWP7T port map(I => TL01_CLR1_n_510, ZN => TL01_CLR1_n_511);
  TL01_CLR1_g41506 : INVD0BWP7T port map(I => TL01_CLR1_n_502, ZN => TL01_CLR1_n_501);
  TL01_CLR1_g41507 : INVD0BWP7T port map(I => TL01_CLR1_n_495, ZN => TL01_CLR1_n_494);
  TL01_CLR1_g41508 : INVD1BWP7T port map(I => TL01_CLR1_n_490, ZN => TL01_CLR1_n_491);
  TL01_CLR1_g41509 : INVD0BWP7T port map(I => TL01_CLR1_n_488, ZN => TL01_CLR1_n_487);
  TL01_CLR1_g41511 : INVD1BWP7T port map(I => TL01_CLR1_n_485, ZN => TL01_CLR1_n_484);
  TL01_CLR1_g41512 : FA1D0BWP7T port map(A => hcountintern(2), B => char1posx(1), CI => TL01_CLR1_n_142, CO => TL01_CLR1_n_517, S => TL01_CLR1_n_519);
  TL01_CLR1_g41513 : FA1D0BWP7T port map(A => hcountintern(2), B => char2posx(1), CI => TL01_CLR1_n_143, CO => TL01_CLR1_n_515, S => TL01_CLR1_n_516);
  TL01_CLR1_g41514 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_359, A2 => TL01_CLR1_n_173, ZN => TL01_CLR1_n_483);
  TL01_CLR1_g41515 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_161, A2 => TL01_CLR1_n_346, B => TL01_CLR1_n_263, ZN => TL01_CLR1_n_482);
  TL01_CLR1_g41516 : AOI211XD0BWP7T port map(A1 => TL01_CLR1_n_195, A2 => TL01_CLR1_n_52, B => char1posy(1), C => char1posy(0), ZN => TL01_CLR1_n_481);
  TL01_CLR1_g41517 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_363, A2 => TL01_CLR1_n_332, ZN => TL01_CLR1_n_480);
  TL01_CLR1_g41518 : AO21D0BWP7T port map(A1 => TL01_CLR1_n_332, A2 => TL01_CLR1_n_1486, B => TL01_CLR1_n_1488, Z => TL01_CLR1_n_479);
  TL01_CLR1_g41519 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_399, A2 => TL01_CLR1_n_415, ZN => TL01_CLR1_n_478);
  TL01_CLR1_g41520 : IND4D0BWP7T port map(A1 => TL01_CLR1_n_121, B1 => char2perc(3), B2 => FE_DBTN6_char2perc_2, B3 => TL01_CLR1_n_224, ZN => TL01_CLR1_n_477);
  TL01_CLR1_g41521 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_293, A2 => TL01_CLR1_n_192, B => TL01_CLR1_n_425, ZN => TL01_CLR1_n_476);
  TL01_CLR1_g41522 : AO21D0BWP7T port map(A1 => TL01_CLR1_n_128, A2 => char2posy(0), B => TL01_CLR1_n_203, Z => TL01_CLR1_n_475);
  TL01_CLR1_g41523 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_304, A2 => TL01_CLR1_n_329, B => TL01_CLR1_n_372, ZN => TL01_CLR1_n_1475);
  TL01_CLR1_g41524 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_302, A2 => TL01_CLR1_n_331, B => TL01_CLR1_n_370, ZN => TL01_CLR1_n_1484);
  TL01_CLR1_g41525 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_405, B1 => TL01_CLR1_n_327, ZN => TL01_CLR1_n_514);
  TL01_CLR1_g41526 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_412, A2 => TL01_CLR1_n_234, ZN => TL01_CLR1_n_513);
  TL01_CLR1_g41527 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_415, B1 => TL01_CLR1_n_395, ZN => TL01_CLR1_n_512);
  TL01_CLR1_g41528 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_375, A2 => TL01_CLR1_n_317, ZN => TL01_CLR1_n_510);
  TL01_CLR1_g41529 : IAO21D0BWP7T port map(A1 => TL01_CLR1_n_118, A2 => FE_DBTN0_char2posx_0, B => char2posx(3), ZN => TL01_CLR1_n_509);
  TL01_CLR1_g41530 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_408, A2 => TL01_CLR1_n_197, Z => TL01_CLR1_n_508);
  TL01_CLR1_g41531 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_258, A2 => hcountintern(3), ZN => TL01_CLR1_n_507);
  TL01_CLR1_g41532 : INR2D1BWP7T port map(A1 => TL01_CLR1_n_382, B1 => TL01_CLR1_n_152, ZN => TL01_CLR1_n_506);
  TL01_CLR1_g41533 : INR2D1BWP7T port map(A1 => TL01_CLR1_n_380, B1 => TL01_CLR1_n_99, ZN => TL01_CLR1_n_505);
  TL01_CLR1_g41534 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_433, A2 => TL01_CLR1_n_190, ZN => TL01_CLR1_n_504);
  TL01_CLR1_g41535 : OAI211D1BWP7T port map(A1 => char2posy(0), A2 => TL01_CLR1_n_57, B => TL01_CLR1_n_272, C => TL01_CLR1_n_159, ZN => TL01_CLR1_n_503);
  TL01_CLR1_g41536 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_374, A2 => TL01_CLR1_n_285, ZN => TL01_CLR1_n_502);
  TL01_CLR1_g41537 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_432, A2 => TL01_CLR1_n_190, ZN => TL01_CLR1_n_500);
  TL01_CLR1_g41538 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_433, A2 => TL01_CLR1_n_349, ZN => TL01_CLR1_n_499);
  TL01_CLR1_g41539 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_399, A2 => TL01_CLR1_n_324, ZN => TL01_CLR1_n_498);
  TL01_CLR1_g41540 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_433, A2 => TL01_CLR1_n_190, ZN => TL01_CLR1_n_497);
  TL01_CLR1_g41541 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_256, A2 => TL01_CLR1_n_54, ZN => TL01_CLR1_n_496);
  TL01_CLR1_g41542 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_414, A2 => TL01_CLR1_n_51, ZN => TL01_CLR1_n_495);
  TL01_CLR1_g41544 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_307, A2 => TL01_CLR1_n_415, ZN => TL01_CLR1_n_493);
  TL01_CLR1_g41545 : AOI21D1BWP7T port map(A1 => TL01_CLR1_n_187, A2 => TL01_CLR1_n_99, B => TL01_CLR1_n_61, ZN => TL01_CLR1_n_492);
  TL01_CLR1_g41546 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_414, A2 => TL01_hcount_int(0), ZN => TL01_CLR1_n_490);
  TL01_CLR1_g41547 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_407, A2 => TL01_CLR1_n_315, ZN => TL01_CLR1_n_489);
  TL01_CLR1_g41548 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_402, A2 => TL01_CLR1_n_51, ZN => TL01_CLR1_n_488);
  TL01_CLR1_g41549 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_402, A2 => TL01_hcount_int(0), Z => TL01_CLR1_n_486);
  TL01_CLR1_g41551 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_393, A2 => vcountintern(3), ZN => TL01_CLR1_n_485);
  TL01_CLR1_g41552 : INVD1BWP7T port map(I => TL01_CLR1_n_468, ZN => TL01_CLR1_n_469);
  TL01_CLR1_g41553 : INVD1BWP7T port map(I => TL01_CLR1_n_456, ZN => TL01_CLR1_n_455);
  TL01_CLR1_g41554 : AOI32D1BWP7T port map(A1 => TL01_CLR1_n_240, A2 => TL01_CLR1_n_175, A3 => TL01_CLR1_n_56, B1 => TL01_CLR1_n_252, B2 => TL01_CLR1_n_110, ZN => TL01_CLR1_n_454);
  TL01_CLR1_g41555 : AO21D0BWP7T port map(A1 => TL01_CLR1_n_328, A2 => TL01_CLR1_n_1477, B => TL01_CLR1_n_1479, Z => TL01_CLR1_n_453);
  TL01_CLR1_g41556 : OA21D0BWP7T port map(A1 => TL01_CLR1_n_1489, A2 => TL01_CLR1_n_95, B => TL01_CLR1_n_370, Z => TL01_CLR1_n_452);
  TL01_CLR1_g41557 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_191, A2 => FE_DBTN10_char1perc_1, B1 => TL01_CLR1_n_342, B2 => TL01_CLR1_n_56, ZN => TL01_CLR1_n_451);
  TL01_CLR1_g41558 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_269, A2 => TL01_CLR1_n_130, B => TL01_CLR1_n_218, ZN => TL01_CLR1_n_450);
  TL01_CLR1_g41559 : OA21D0BWP7T port map(A1 => TL01_CLR1_n_1480, A2 => TL01_CLR1_n_73, B => TL01_CLR1_n_372, Z => TL01_CLR1_n_449);
  TL01_CLR1_g41560 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_108, A2 => TL01_CLR1_n_133, B1 => TL01_CLR1_n_250, B2 => char1perc(1), ZN => TL01_CLR1_n_448);
  TL01_CLR1_g41561 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_195, A2 => TL01_CLR1_n_351, B => TL01_CLR1_n_52, ZN => TL01_CLR1_n_447);
  TL01_CLR1_g41562 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_351, A2 => char1posy(0), B => TL01_CLR1_n_195, ZN => TL01_CLR1_n_446);
  TL01_CLR1_g41563 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_300, A2 => TL01_CLR1_n_102, B => TL01_CLR1_n_426, ZN => TL01_CLR1_n_445);
  TL01_CLR1_g41564 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_292, A2 => TL01_CLR1_n_340, B => TL01_CLR1_n_299, ZN => TL01_CLR1_n_444);
  TL01_CLR1_g41565 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_250, A2 => TL01_CLR1_n_155, B1 => TL01_CLR1_n_301, B2 => TL01_CLR1_n_191, ZN => TL01_CLR1_n_443);
  TL01_CLR1_g41566 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_273, A2 => FE_DBTN13_char1perc_5, B1 => TL01_CLR1_n_119, B2 => char1perc(5), ZN => TL01_CLR1_n_442);
  TL01_CLR1_g41567 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_133, A2 => char1perc(3), B1 => TL01_CLR1_n_151, B2 => char1perc(1), ZN => TL01_CLR1_n_441);
  TL01_CLR1_g41568 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_184, A2 => TL01_CLR1_n_65, B => TL01_CLR1_n_159, ZN => TL01_CLR1_n_440);
  TL01_CLR1_g41569 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_270, A2 => hcountintern(9), B1 => TL01_CLR1_n_150, B2 => TL01_CLR1_n_123, ZN => TL01_CLR1_n_439);
  TL01_CLR1_g41570 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_229, A2 => TL01_CLR1_n_120, B1 => TL01_CLR1_n_136, B2 => TL01_CLR1_n_99, ZN => TL01_CLR1_n_438);
  TL01_CLR1_g41571 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_134, A2 => char2perc(3), B1 => TL01_CLR1_n_345, B2 => char2perc(1), ZN => TL01_CLR1_n_437);
  TL01_CLR1_g41572 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_333, A2 => vcountintern(3), B1 => TL01_CLR1_n_176, B2 => TL01_CLR1_n_52, ZN => TL01_CLR1_n_436);
  TL01_CLR1_g41573 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_277, A2 => char1perc(5), B1 => TL01_CLR1_n_223, B2 => TL01_CLR1_n_131, ZN => TL01_CLR1_n_435);
  TL01_CLR1_g41574 : IND3D1BWP7T port map(A1 => inputsp2(2), B1 => TL01_CLR1_n_202, B2 => TL01_CLR1_n_372, ZN => TL01_CLR1_n_474);
  TL01_CLR1_g41575 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_341, A2 => vcountintern(3), B => TL01_CLR1_n_416, ZN => TL01_CLR1_n_473);
  TL01_CLR1_g41576 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_431, A2 => TL01_CLR1_n_159, ZN => TL01_CLR1_n_434);
  TL01_CLR1_g41577 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_301, A2 => TL01_CLR1_n_156, B1 => TL01_CLR1_n_292, B2 => TL01_CLR1_n_151, ZN => TL01_CLR1_n_472);
  TL01_CLR1_g41578 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_343, A2 => TL01_CLR1_n_346, B1 => TL01_CLR1_n_347, B2 => TL01_CLR1_n_172, ZN => TL01_CLR1_n_471);
  TL01_CLR1_g41579 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_201, A2 => TL01_CLR1_n_191, B1 => TL01_CLR1_n_152, B2 => TL01_CLR1_n_171, ZN => TL01_CLR1_n_470);
  TL01_CLR1_g41580 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_196, A2 => TL01_CLR1_n_347, B1 => TL01_CLR1_n_172, B2 => TL01_CLR1_n_99, ZN => TL01_CLR1_n_468);
  TL01_CLR1_g41581 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_204, A2 => TL01_CLR1_n_52, B1 => TL01_CLR1_n_204, B2 => TL01_CLR1_n_52, ZN => TL01_CLR1_n_467);
  TL01_CLR1_g41582 : IND3D1BWP7T port map(A1 => inputsp1(2), B1 => TL01_CLR1_n_207, B2 => TL01_CLR1_n_370, ZN => TL01_CLR1_n_466);
  TL01_CLR1_g41583 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_1562, A2 => TL01_CLR1_n_52, B1 => TL01_CLR1_n_1562, B2 => TL01_CLR1_n_52, ZN => TL01_CLR1_n_465);
  TL01_CLR1_g41584 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_181, A2 => char2posx(2), B1 => TL01_CLR1_n_181, B2 => char2posx(2), ZN => TL01_CLR1_n_464);
  TL01_CLR1_g41585 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_137, A2 => char1posx(2), B1 => TL01_CLR1_n_137, B2 => char1posx(2), ZN => TL01_CLR1_n_463);
  TL01_CLR1_g41586 : IAO21D0BWP7T port map(A1 => TL01_CLR1_n_177, A2 => TL01_CLR1_n_69, B => char1posx(3), ZN => TL01_CLR1_n_462);
  TL01_CLR1_g41587 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_118, A2 => char2posx(3), B1 => TL01_CLR1_n_118, B2 => char2posx(3), ZN => TL01_CLR1_n_461);
  TL01_CLR1_g41588 : AOI32D1BWP7T port map(A1 => TL01_CLR1_n_104, A2 => TL01_CLR1_n_146, A3 => hcountintern(4), B1 => TL01_CLR1_n_281, B2 => TL01_CLR1_n_53, ZN => TL01_CLR1_n_460);
  TL01_CLR1_g41589 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_177, A2 => char1posx(3), B1 => TL01_CLR1_n_177, B2 => char1posx(3), ZN => TL01_CLR1_n_459);
  TL01_CLR1_g41590 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_125, A2 => FE_DBTN2_char1posy_3, B => TL01_CLR1_n_420, ZN => TL01_CLR1_n_458);
  TL01_CLR1_g41591 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_128, A2 => char2posy(3), B => TL01_CLR1_n_417, ZN => TL01_CLR1_n_457);
  TL01_CLR1_g41592 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_217, A2 => TL01_CLR1_n_141, B1 => TL01_CLR1_n_217, B2 => TL01_CLR1_n_141, ZN => TL01_CLR1_n_456);
  TL01_CLR1_g41593 : INVD1BWP7T port map(I => TL01_CLR1_n_433, ZN => TL01_CLR1_n_432);
  TL01_CLR1_g41594 : INVD0BWP7T port map(I => TL01_CLR1_n_426, ZN => TL01_CLR1_n_427);
  TL01_CLR1_g41595 : INVD0BWP7T port map(I => TL01_CLR1_n_417, ZN => TL01_CLR1_n_418);
  TL01_CLR1_g41596 : INVD0BWP7T port map(I => TL01_CLR1_n_412, ZN => TL01_CLR1_n_411);
  TL01_CLR1_g41597 : INVD0BWP7T port map(I => TL01_CLR1_n_410, ZN => TL01_CLR1_n_409);
  TL01_CLR1_g41598 : INVD0BWP7T port map(I => TL01_CLR1_n_407, ZN => TL01_CLR1_n_406);
  TL01_CLR1_g41599 : INVD0BWP7T port map(I => TL01_CLR1_n_404, ZN => TL01_CLR1_n_403);
  TL01_CLR1_g41600 : INVD0BWP7T port map(I => TL01_CLR1_n_401, ZN => TL01_CLR1_n_400);
  TL01_CLR1_g41601 : INVD0BWP7T port map(I => TL01_CLR1_n_399, ZN => TL01_CLR1_n_398);
  TL01_CLR1_g41602 : INVD1BWP7T port map(I => TL01_CLR1_n_397, ZN => TL01_CLR1_n_396);
  TL01_CLR1_g41603 : INVD1BWP7T port map(I => TL01_CLR1_n_395, ZN => TL01_CLR1_n_394);
  TL01_CLR1_g41604 : HA1D0BWP7T port map(A => TL01_CLR1_n_57, B => TL01_CLR1_n_115, CO => TL01_CLR1_n_393, S => TL01_CLR1_n_433);
  TL01_CLR1_g41605 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_295, A2 => TL01_CLR1_n_1494, ZN => TL01_CLR1_n_392);
  TL01_CLR1_g41606 : ND2D0BWP7T port map(A1 => TL01_CLR1_n_102, A2 => TL01_CLR1_n_138, ZN => TL01_CLR1_n_391);
  TL01_CLR1_g41607 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_184, B1 => char1posy(1), ZN => TL01_CLR1_n_431);
  TL01_CLR1_g41608 : NR2D0BWP7T port map(A1 => TL01_CLR1_n_307, A2 => TL01_CLR1_n_246, ZN => TL01_CLR1_n_430);
  TL01_CLR1_g41609 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_337, A2 => TL01_CLR1_n_260, ZN => TL01_CLR1_n_429);
  TL01_CLR1_g41610 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_110, A2 => TL01_CLR1_n_178, ZN => TL01_CLR1_n_428);
  TL01_CLR1_g41611 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_293, A2 => TL01_CLR1_n_345, ZN => TL01_CLR1_n_426);
  TL01_CLR1_g41612 : NR2D0BWP7T port map(A1 => TL01_CLR1_n_242, A2 => TL01_CLR1_n_102, ZN => TL01_CLR1_n_425);
  TL01_CLR1_g41613 : INR2XD0BWP7T port map(A1 => char2posx(3), B1 => TL01_CLR1_n_118, ZN => TL01_CLR1_n_424);
  TL01_CLR1_g41614 : INR2D1BWP7T port map(A1 => char1posx(3), B1 => TL01_CLR1_n_177, ZN => TL01_CLR1_n_423);
  TL01_CLR1_g41615 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_163, A2 => TL01_CLR1_n_99, ZN => TL01_CLR1_n_422);
  TL01_CLR1_g41616 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_240, A2 => TL01_CLR1_n_340, ZN => TL01_CLR1_n_421);
  TL01_CLR1_g41617 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_125, A2 => FE_DBTN2_char1posy_3, ZN => TL01_CLR1_n_420);
  TL01_CLR1_g41618 : NR2D0BWP7T port map(A1 => TL01_CLR1_n_172, A2 => TL01_CLR1_n_102, ZN => TL01_CLR1_n_419);
  TL01_CLR1_g41619 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_128, A2 => char2posy(3), ZN => TL01_CLR1_n_417);
  TL01_CLR1_g41621 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_341, A2 => vcountintern(3), ZN => TL01_CLR1_n_416);
  TL01_CLR1_g41622 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_319, A2 => TL01_CLR1_n_238, ZN => TL01_CLR1_n_415);
  TL01_CLR1_g41624 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_317, A2 => hcountintern(4), ZN => TL01_CLR1_n_414);
  TL01_CLR1_g41625 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_324, A2 => TL01_hcount_int(0), ZN => TL01_CLR1_n_413);
  TL01_CLR1_g41626 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_309, A2 => TL01_hcount_int(0), ZN => TL01_CLR1_n_412);
  TL01_CLR1_g41627 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_230, A2 => TL01_CLR1_n_152, B => TL01_CLR1_n_87, ZN => TL01_CLR1_n_410);
  TL01_CLR1_g41628 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_313, A2 => hcountintern(4), ZN => TL01_CLR1_n_408);
  TL01_CLR1_g41629 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_325, A2 => TL01_hcount_int(0), ZN => TL01_CLR1_n_407);
  TL01_CLR1_g41630 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_286, A2 => hcountintern(4), ZN => TL01_CLR1_n_405);
  TL01_CLR1_g41631 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_317, A2 => TL01_hcount_int(0), ZN => TL01_CLR1_n_404);
  TL01_CLR1_g41632 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_308, A2 => TL01_CLR1_n_53, ZN => TL01_CLR1_n_402);
  TL01_CLR1_g41633 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_330, A2 => TL01_hcount_int(0), ZN => TL01_CLR1_n_401);
  TL01_CLR1_g41634 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_290, A2 => TL01_hcount_int(0), ZN => TL01_CLR1_n_399);
  TL01_CLR1_g41635 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_327, A2 => TL01_CLR1_n_337, ZN => TL01_CLR1_n_397);
  TL01_CLR1_g41636 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_330, A2 => TL01_CLR1_n_51, ZN => TL01_CLR1_n_395);
  TL01_CLR1_g41637 : INVD0BWP7T port map(I => TL01_CLR1_n_388, ZN => TL01_CLR1_n_389);
  TL01_CLR1_g41638 : INVD1BWP7T port map(I => TL01_CLR1_n_377, ZN => TL01_CLR1_n_376);
  TL01_CLR1_g41639 : INVD0BWP7T port map(I => TL01_CLR1_n_374, ZN => TL01_CLR1_n_373);
  TL01_CLR1_g41640 : INVD0BWP7T port map(I => TL01_CLR1_n_372, ZN => TL01_CLR1_n_371);
  TL01_CLR1_g41641 : INVD0BWP7T port map(I => TL01_CLR1_n_370, ZN => TL01_CLR1_n_369);
  TL01_CLR1_g41642 : INVD0BWP7T port map(I => TL01_CLR1_n_368, ZN => TL01_CLR1_n_367);
  TL01_CLR1_g41643 : NR3D0BWP7T port map(A1 => TL01_CLR1_n_249, A2 => TL01_CLR1_n_52, A3 => TL01_CLR1_n_83, ZN => TL01_CLR1_n_366);
  TL01_CLR1_g41644 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_216, A2 => FE_DBTN11_char1perc_3, B1 => TL01_CLR1_n_179, B2 => TL01_CLR1_n_182, ZN => TL01_CLR1_n_365);
  TL01_CLR1_g41645 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_255, A2 => TL01_CLR1_n_100, B1 => TL01_CLR1_n_255, B2 => TL01_CLR1_n_124, ZN => TL01_CLR1_n_364);
  TL01_CLR1_g41646 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_208, A2 => TL01_CLR1_char1_sprite_frame_control_state_2, B1 => TL01_CLR1_n_97, B2 => FE_PHN106_TL01_CLR1_char1_sprite_frame_control_state_0, ZN => TL01_CLR1_n_363);
  TL01_CLR1_g41647 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_202, A2 => TL01_CLR1_n_117, B1 => TL01_CLR1_n_135, B2 => inputsp2(3), ZN => TL01_CLR1_n_362);
  TL01_CLR1_g41648 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_231, A2 => hcountintern(7), B1 => TL01_CLR1_n_220, B2 => TL01_CLR1_n_82, ZN => TL01_CLR1_n_361);
  TL01_CLR1_g41649 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_264, A2 => TL01_CLR1_n_130, B => TL01_CLR1_n_179, ZN => TL01_CLR1_n_360);
  TL01_CLR1_g41650 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_221, A2 => TL01_CLR1_n_161, B => TL01_CLR1_n_140, ZN => TL01_CLR1_n_359);
  TL01_CLR1_g41651 : NR4D0BWP7T port map(A1 => TL01_CLR1_n_132, A2 => FE_DBTN13_char1perc_5, A3 => char1perc(7), A4 => char1perc(6), ZN => TL01_CLR1_n_358);
  TL01_CLR1_g41652 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_262, A2 => TL01_CLR1_n_154, A3 => TL01_CLR1_n_100, ZN => TL01_CLR1_n_357);
  TL01_CLR1_g41653 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_219, A2 => TL01_CLR1_n_154, B => hcountintern(7), ZN => TL01_CLR1_n_356);
  TL01_CLR1_g41654 : IND3D1BWP7T port map(A1 => TL01_CLR1_n_119, B1 => char1perc(3), B2 => TL01_CLR1_n_222, ZN => TL01_CLR1_n_355);
  TL01_CLR1_g41655 : OAI211D1BWP7T port map(A1 => char1perc(5), A2 => TL01_CLR1_n_109, B => FE_DBTN12_char1perc_4, C => char1perc(7), ZN => TL01_CLR1_n_354);
  TL01_CLR1_g41656 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_224, A2 => TL01_CLR1_n_77, B => TL01_CLR1_n_99, ZN => TL01_CLR1_n_353);
  TL01_CLR1_g41657 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_77, A2 => FE_DBTN6_char2perc_2, B => TL01_CLR1_n_99, ZN => TL01_CLR1_n_352);
  TL01_CLR1_g41658 : AO211D0BWP7T port map(A1 => FE_DBTN9_char2perc_5, A2 => char2perc(6), B => TL01_CLR1_n_120, C => FE_DBTN8_char2perc_4, Z => TL01_CLR1_n_390);
  TL01_CLR1_g41659 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_285, A2 => TL01_CLR1_n_232, ZN => TL01_CLR1_n_388);
  TL01_CLR1_g41660 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_283, A2 => TL01_CLR1_n_238, ZN => TL01_CLR1_n_387);
  TL01_CLR1_g41661 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_195, A2 => char1posy(3), B1 => TL01_CLR1_n_195, B2 => char1posy(3), ZN => TL01_CLR1_n_386);
  TL01_CLR1_g41662 : CKAN2D1BWP7T port map(A1 => TL01_CLR1_n_290, A2 => TL01_CLR1_n_284, Z => TL01_CLR1_n_385);
  TL01_CLR1_g41663 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_203, A2 => char2posy(3), B1 => TL01_CLR1_n_203, B2 => char2posy(3), ZN => TL01_CLR1_n_384);
  TL01_CLR1_g41664 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_226, A2 => char1perc(4), B1 => TL01_CLR1_n_164, B2 => FE_DBTN12_char1perc_4, ZN => TL01_CLR1_n_383);
  TL01_CLR1_g41665 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_226, A2 => FE_DBTN12_char1perc_4, B1 => TL01_CLR1_n_108, B2 => char1perc(4), ZN => TL01_CLR1_n_382);
  TL01_CLR1_g41666 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_225, A2 => char2perc(4), B1 => TL01_CLR1_n_163, B2 => FE_DBTN8_char2perc_4, ZN => TL01_CLR1_n_381);
  TL01_CLR1_g41667 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_225, A2 => FE_DBTN8_char2perc_4, B1 => TL01_CLR1_n_161, B2 => char2perc(4), ZN => TL01_CLR1_n_380);
  TL01_CLR1_g41668 : CKND2D1BWP7T port map(A1 => TL01_CLR1_n_311, A2 => TL01_CLR1_n_314, ZN => TL01_CLR1_n_379);
  TL01_CLR1_g41669 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_215, A2 => TL01_CLR1_n_180, B1 => TL01_CLR1_n_215, B2 => TL01_CLR1_n_180, ZN => TL01_CLR1_n_378);
  TL01_CLR1_g41670 : CKND2D1BWP7T port map(A1 => TL01_CLR1_n_313, A2 => TL01_CLR1_n_306, ZN => TL01_CLR1_n_377);
  TL01_CLR1_g41671 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_308, A2 => TL01_hcount_int(0), ZN => TL01_CLR1_n_375);
  TL01_CLR1_g41672 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_322, A2 => TL01_CLR1_n_319, ZN => TL01_CLR1_n_374);
  TL01_CLR1_g41673 : INR4D0BWP7T port map(A1 => TL01_CLR1_n_1478, B1 => TL01_CLR1_char2_sprite_frame_control_frame_count_4, B2 => TL01_CLR1_char2_sprite_frame_control_frame_count_3, B3 => TL01_CLR1_char2_sprite_frame_control_frame_count_2, ZN => TL01_CLR1_n_372);
  TL01_CLR1_g41674 : INR4D0BWP7T port map(A1 => TL01_CLR1_n_1487, B1 => TL01_CLR1_char1_sprite_frame_control_frame_count_4, B2 => FE_PHN109_TL01_CLR1_char1_sprite_frame_control_frame_count_3, B3 => FE_PHN111_TL01_CLR1_char1_sprite_frame_control_frame_count_2, ZN => TL01_CLR1_n_370);
  TL01_CLR1_g41675 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_285, A2 => TL01_CLR1_n_286, ZN => TL01_CLR1_n_368);
  TL01_CLR1_g41676 : INVD0BWP7T port map(I => TL01_CLR1_n_125, ZN => TL01_CLR1_n_351);
  TL01_CLR1_g41677 : INVD0BWP7T port map(I => TL01_CLR1_n_212, ZN => TL01_CLR1_n_350);
  TL01_CLR1_g41678 : INVD1BWP7T port map(I => TL01_CLR1_n_190, ZN => TL01_CLR1_n_349);
  TL01_CLR1_g41679 : INVD0BWP7T port map(I => TL01_CLR1_n_116, ZN => TL01_CLR1_n_348);
  TL01_CLR1_g41680 : INVD1BWP7T port map(I => TL01_CLR1_n_192, ZN => TL01_CLR1_n_347);
  TL01_CLR1_g41681 : INVD0BWP7T port map(I => TL01_CLR1_n_102, ZN => TL01_CLR1_n_346);
  TL01_CLR1_g41682 : INVD1BWP7T port map(I => TL01_CLR1_n_99, ZN => TL01_CLR1_n_345);
  TL01_CLR1_g41684 : INVD1BWP7T port map(I => TL01_CLR1_n_196, ZN => TL01_CLR1_n_343);
  TL01_CLR1_g41685 : INVD1BWP7T port map(I => TL01_CLR1_n_201, ZN => TL01_CLR1_n_342);
  TL01_CLR1_g41686 : INVD0BWP7T port map(I => TL01_CLR1_n_159, ZN => TL01_CLR1_n_341);
  TL01_CLR1_g41687 : INVD0BWP7T port map(I => TL01_CLR1_n_191, ZN => TL01_CLR1_n_340);
  TL01_CLR1_g41690 : INVD0BWP7T port map(I => TL01_CLR1_n_331, ZN => TL01_CLR1_n_332);
  TL01_CLR1_g41691 : INVD0BWP7T port map(I => TL01_CLR1_n_329, ZN => TL01_CLR1_n_328);
  TL01_CLR1_g41692 : INVD1BWP7T port map(I => TL01_CLR1_n_325, ZN => TL01_CLR1_n_324);
  TL01_CLR1_g41693 : INVD0BWP7T port map(I => TL01_CLR1_n_323, ZN => TL01_CLR1_n_322);
  TL01_CLR1_g41694 : INVD1BWP7T port map(I => TL01_CLR1_n_321, ZN => TL01_CLR1_n_320);
  TL01_CLR1_g41695 : INVD0BWP7T port map(I => TL01_CLR1_n_319, ZN => TL01_CLR1_n_318);
  TL01_CLR1_g41696 : INVD1BWP7T port map(I => TL01_CLR1_n_317, ZN => TL01_CLR1_n_316);
  TL01_CLR1_g41697 : INVD1BWP7T port map(I => TL01_CLR1_n_315, ZN => TL01_CLR1_n_314);
  TL01_CLR1_g41698 : INVD0BWP7T port map(I => TL01_CLR1_n_313, ZN => TL01_CLR1_n_312);
  TL01_CLR1_g41699 : INVD1BWP7T port map(I => TL01_CLR1_n_311, ZN => TL01_CLR1_n_310);
  TL01_CLR1_g41700 : INVD1BWP7T port map(I => TL01_CLR1_n_309, ZN => TL01_CLR1_n_308);
  TL01_CLR1_g41701 : INVD1BWP7T port map(I => TL01_CLR1_n_307, ZN => TL01_CLR1_n_306);
  TL01_CLR1_g41702 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_1488, A2 => TL01_CLR1_n_261, ZN => FE_PHN149_TL01_CLR1_n_305);
  TL01_CLR1_g41703 : INR2D1BWP7T port map(A1 => TL01_CLR1_n_202, B1 => inputsp2(3), ZN => TL01_CLR1_n_304);
  TL01_CLR1_g41704 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_268, A2 => TL01_CLR1_n_1479, ZN => TL01_CLR1_n_303);
  TL01_CLR1_g41705 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_208, A2 => inputsp1(3), ZN => TL01_CLR1_n_302);
  TL01_CLR1_g41706 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_202, A2 => inputsp2(2), ZN => TL01_CLR1_n_339);
  TL01_CLR1_g41707 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_207, A2 => inputsp1(2), ZN => TL01_CLR1_n_338);
  TL01_CLR1_g41708 : IND2D1BWP7T port map(A1 => TL01_CLR1_char1_sprite_frame_control_frame_count_4, B1 => TL01_CLR1_n_186, ZN => TL01_CLR1_n_1486);
  TL01_CLR1_g41709 : CKAN2D1BWP7T port map(A1 => TL01_CLR1_n_249, A2 => vcountintern(3), Z => TL01_CLR1_n_337);
  TL01_CLR1_g41710 : IND2D1BWP7T port map(A1 => TL01_CLR1_char2_sprite_frame_control_frame_count_4, B1 => TL01_CLR1_n_189, ZN => TL01_CLR1_n_1477);
  TL01_CLR1_g41711 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_195, A2 => FE_DBTN2_char1posy_3, Z => TL01_CLR1_n_336);
  TL01_CLR1_g41712 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_203, B1 => char2posy(3), ZN => TL01_CLR1_n_335);
  TL01_CLR1_g41713 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_247, A2 => TL01_hcount_int(0), ZN => TL01_CLR1_n_334);
  TL01_CLR1_g41714 : CKAN2D1BWP7T port map(A1 => TL01_CLR1_n_249, A2 => TL01_CLR1_n_83, Z => TL01_CLR1_n_333);
  TL01_CLR1_g41715 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_214, A2 => TL01_CLR1_n_95, ZN => TL01_CLR1_n_331);
  TL01_CLR1_g41716 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_235, A2 => hcountintern(4), ZN => TL01_CLR1_n_330);
  TL01_CLR1_g41717 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_213, A2 => TL01_CLR1_n_73, ZN => TL01_CLR1_n_329);
  TL01_CLR1_g41718 : IND2D1BWP7T port map(A1 => inputsp2(3), B1 => TL01_CLR1_n_213, ZN => TL01_CLR1_n_1480);
  TL01_CLR1_g41719 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_214, A2 => TL01_CLR1_n_97, ZN => TL01_CLR1_n_1489);
  TL01_CLR1_g41720 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_249, A2 => vcountintern(3), ZN => TL01_CLR1_n_327);
  TL01_CLR1_g41721 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_255, A2 => hcountintern(4), ZN => TL01_CLR1_n_326);
  TL01_CLR1_g41722 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_248, A2 => hcountintern(4), ZN => TL01_CLR1_n_325);
  TL01_CLR1_g41723 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_238, A2 => TL01_hcount_int(0), ZN => TL01_CLR1_n_323);
  TL01_CLR1_g41724 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_253, A2 => TL01_CLR1_n_104, ZN => TL01_CLR1_n_321);
  TL01_CLR1_g41725 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_236, A2 => TL01_hcount_int(0), ZN => TL01_CLR1_n_319);
  TL01_CLR1_g41726 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_254, A2 => hcountintern(1), ZN => TL01_CLR1_n_317);
  TL01_CLR1_g41727 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_247, A2 => TL01_CLR1_n_51, ZN => TL01_CLR1_n_315);
  TL01_CLR1_g41728 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_246, A2 => TL01_hcount_int(0), ZN => TL01_CLR1_n_313);
  TL01_CLR1_g41729 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_232, A2 => TL01_CLR1_n_51, ZN => TL01_CLR1_n_311);
  TL01_CLR1_g41730 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_254, A2 => TL01_CLR1_n_85, ZN => TL01_CLR1_n_309);
  TL01_CLR1_g41731 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_235, A2 => TL01_hcount_int(0), ZN => TL01_CLR1_n_307);
  TL01_CLR1_g41732 : INVD0BWP7T port map(I => TL01_CLR1_n_295, ZN => TL01_CLR1_n_294);
  TL01_CLR1_g41733 : INVD0BWP7T port map(I => TL01_CLR1_n_288, ZN => TL01_CLR1_n_287);
  TL01_CLR1_g41734 : INVD0BWP7T port map(I => TL01_CLR1_n_285, ZN => TL01_CLR1_n_284);
  TL01_CLR1_g41736 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_101, A2 => hcountintern(8), B => TL01_CLR1_n_153, ZN => TL01_CLR1_n_282);
  TL01_CLR1_g41737 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_104, A2 => TL01_CLR1_n_54, B => TL01_CLR1_n_146, ZN => TL01_CLR1_n_281);
  TL01_CLR1_g41738 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_149, A2 => hcountintern(4), B => TL01_CLR1_n_157, ZN => TL01_CLR1_n_280);
  TL01_CLR1_g41739 : IOA21D1BWP7T port map(A1 => inputsp2(2), A2 => inputsp2(3), B => TL01_CLR1_n_213, ZN => TL01_CLR1_n_279);
  TL01_CLR1_g41740 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_95, A2 => TL01_CLR1_n_97, B => TL01_CLR1_n_214, ZN => TL01_CLR1_n_278);
  TL01_CLR1_g41741 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_119, A2 => TL01_CLR1_n_132, B => TL01_CLR1_n_266, ZN => TL01_CLR1_n_277);
  TL01_CLR1_g41742 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_129, A2 => TL01_CLR1_n_155, A3 => char1perc(5), ZN => TL01_CLR1_n_276);
  TL01_CLR1_g41743 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_121, A2 => TL01_CLR1_n_173, B => TL01_CLR1_n_263, ZN => TL01_CLR1_n_275);
  TL01_CLR1_g41744 : AO21D0BWP7T port map(A1 => TL01_CLR1_n_109, A2 => TL01_CLR1_n_156, B => TL01_CLR1_n_265, Z => TL01_CLR1_n_274);
  TL01_CLR1_g41745 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_131, A2 => char1perc(2), B => TL01_CLR1_n_267, ZN => TL01_CLR1_n_273);
  TL01_CLR1_g41746 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_180, A2 => vcountintern(2), B => char2posy(1), ZN => TL01_CLR1_n_272);
  TL01_CLR1_g41747 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_168, A2 => hcountintern(6), B => hcountintern(7), ZN => TL01_CLR1_n_271);
  TL01_CLR1_g41748 : NR3D0BWP7T port map(A1 => TL01_CLR1_n_150, A2 => TL01_CLR1_n_158, A3 => TL01_CLR1_n_100, ZN => TL01_CLR1_n_270);
  TL01_CLR1_g41749 : MOAI22D0BWP7T port map(A1 => FE_DBTN13_char1perc_5, A2 => TL01_CLR1_n_56, B1 => TL01_CLR1_n_151, B2 => char1perc(2), ZN => TL01_CLR1_n_269);
  TL01_CLR1_g41750 : AOI211XD0BWP7T port map(A1 => char1perc(4), A2 => char1perc(2), B => TL01_CLR1_n_130, C => TL01_CLR1_n_129, ZN => TL01_CLR1_n_301);
  TL01_CLR1_g41751 : OA221D0BWP7T port map(A1 => char2perc(4), A2 => char2perc(6), B1 => FE_DBTN6_char2perc_2, B2 => FE_DBTN8_char2perc_4, C => TL01_CLR1_n_127, Z => TL01_CLR1_n_300);
  TL01_CLR1_g41752 : NR2D0BWP7T port map(A1 => TL01_CLR1_n_239, A2 => TL01_CLR1_n_156, ZN => TL01_CLR1_n_299);
  TL01_CLR1_g41753 : NR3D0BWP7T port map(A1 => TL01_CLR1_n_111, A2 => TL01_CLR1_n_164, A3 => char1perc(1), ZN => TL01_CLR1_n_298);
  TL01_CLR1_g41754 : IND3D1BWP7T port map(A1 => TL01_CLR1_n_163, B1 => FE_DBTN5_char2perc_1, B2 => TL01_CLR1_n_112, ZN => TL01_CLR1_n_297);
  TL01_CLR1_g41755 : ND3D0BWP7T port map(A1 => TL01_CLR1_n_112, A2 => char2perc(7), A3 => FE_DBTN7_char2perc_3, ZN => TL01_CLR1_n_296);
  TL01_CLR1_g41756 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_260, A2 => vcountintern(3), ZN => TL01_CLR1_n_295);
  TL01_CLR1_g41757 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_163, A2 => char2perc(4), B => TL01_CLR1_n_162, ZN => TL01_CLR1_n_293);
  TL01_CLR1_g41758 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_164, A2 => char1perc(4), B => TL01_CLR1_n_109, ZN => TL01_CLR1_n_292);
  TL01_CLR1_g41759 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_113, A2 => hcountintern(2), B1 => TL01_CLR1_n_113, B2 => hcountintern(2), ZN => TL01_CLR1_n_291);
  TL01_CLR1_g41760 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_232, A2 => hcountintern(4), ZN => TL01_CLR1_n_290);
  TL01_CLR1_g41761 : AO21D0BWP7T port map(A1 => TL01_CLR1_n_105, A2 => hcountintern(2), B => TL01_CLR1_n_258, Z => TL01_CLR1_n_289);
  TL01_CLR1_g41762 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_234, A2 => TL01_hcount_int(0), ZN => TL01_CLR1_n_288);
  TL01_CLR1_g41763 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_233, A2 => TL01_CLR1_n_51, ZN => TL01_CLR1_n_286);
  TL01_CLR1_g41764 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_237, A2 => TL01_hcount_int(0), ZN => TL01_CLR1_n_285);
  TL01_CLR1_g41765 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_194, A2 => TL01_CLR1_n_197, ZN => TL01_CLR1_n_283);
  TL01_CLR1_g41766 : INVD0BWP7T port map(I => TL01_CLR1_n_265, ZN => TL01_CLR1_n_266);
  TL01_CLR1_g41768 : INVD0BWP7T port map(I => TL01_CLR1_n_254, ZN => TL01_CLR1_n_253);
  TL01_CLR1_g41769 : INVD1BWP7T port map(I => TL01_CLR1_n_248, ZN => TL01_CLR1_n_247);
  TL01_CLR1_g41770 : INVD0BWP7T port map(I => TL01_CLR1_n_246, ZN => TL01_CLR1_n_245);
  TL01_CLR1_g41771 : INVD0BWP7T port map(I => TL01_CLR1_n_1483, ZN => TL01_CLR1_n_2);
  TL01_CLR1_g41772 : INVD0BWP7T port map(I => TL01_CLR1_n_1492, ZN => TL01_CLR1_n_3);
  TL01_CLR1_g41773 : INVD0BWP7T port map(I => TL01_CLR1_n_242, ZN => TL01_CLR1_n_241);
  TL01_CLR1_g41774 : INVD0BWP7T port map(I => TL01_CLR1_n_240, ZN => TL01_CLR1_n_239);
  TL01_CLR1_g41775 : INVD1BWP7T port map(I => TL01_CLR1_n_237, ZN => TL01_CLR1_n_236);
  TL01_CLR1_g41776 : INVD1BWP7T port map(I => TL01_CLR1_n_235, ZN => TL01_CLR1_n_234);
  TL01_CLR1_g41777 : INVD1BWP7T port map(I => TL01_CLR1_n_233, ZN => TL01_CLR1_n_232);
  TL01_CLR1_g41778 : ND2D0BWP7T port map(A1 => TL01_CLR1_n_167, A2 => TL01_CLR1_n_146, ZN => TL01_CLR1_n_231);
  TL01_CLR1_g41779 : ND2D0BWP7T port map(A1 => TL01_CLR1_n_111, A2 => char1perc(7), ZN => TL01_CLR1_n_230);
  TL01_CLR1_g41780 : ND2D0BWP7T port map(A1 => TL01_CLR1_n_173, A2 => TL01_CLR1_n_77, ZN => TL01_CLR1_n_229);
  TL01_CLR1_g41781 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_179, A2 => TL01_CLR1_n_155, Z => TL01_CLR1_n_228);
  TL01_CLR1_g41782 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_117, A2 => TL01_CLR1_char2_sprite_frame_control_state_0, ZN => TL01_CLR1_n_268);
  TL01_CLR1_g41783 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_152, A2 => char1perc(6), ZN => TL01_CLR1_n_267);
  TL01_CLR1_g41784 : NR2D0BWP7T port map(A1 => TL01_CLR1_n_164, A2 => char1perc(7), ZN => TL01_CLR1_n_265);
  TL01_CLR1_g41785 : NR2D0BWP7T port map(A1 => TL01_CLR1_n_108, A2 => TL01_CLR1_n_56, ZN => TL01_CLR1_n_264);
  TL01_CLR1_g41786 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_163, A2 => char2perc(7), Z => TL01_CLR1_n_263);
  TL01_CLR1_g41787 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_145, A2 => hcountintern(5), ZN => TL01_CLR1_n_262);
  TL01_CLR1_g41788 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_1490, B1 => FE_PHN106_TL01_CLR1_char1_sprite_frame_control_state_0, ZN => TL01_CLR1_n_261);
  TL01_CLR1_g41789 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_114, A2 => TL01_CLR1_n_57, ZN => TL01_CLR1_n_260);
  TL01_CLR1_g41790 : IND2D1BWP7T port map(A1 => FE_PHN106_TL01_CLR1_char1_sprite_frame_control_state_0, B1 => TL01_CLR1_n_139, ZN => TL01_CLR1_n_1488);
  TL01_CLR1_g41791 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_1491, B1 => TL01_CLR1_char1_sprite_frame_control_state_2, ZN => TL01_CLR1_n_259);
  TL01_CLR1_g41792 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_105, A2 => hcountintern(2), ZN => TL01_CLR1_n_258);
  TL01_CLR1_g41793 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_135, A2 => FE_PHN99_TL01_CLR1_char2_sprite_frame_control_state_2, ZN => TL01_CLR1_n_257);
  TL01_CLR1_g41794 : IND2D1BWP7T port map(A1 => TL01_CLR1_char2_sprite_frame_control_state_0, B1 => TL01_CLR1_n_185, ZN => TL01_CLR1_n_1479);
  TL01_CLR1_g41795 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_113, B1 => hcountintern(2), ZN => TL01_CLR1_n_256);
  TL01_CLR1_g41796 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_146, A2 => TL01_CLR1_n_113, ZN => TL01_CLR1_n_255);
  TL01_CLR1_g41797 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_150, A2 => hcountintern(2), ZN => TL01_CLR1_n_254);
  TL01_CLR1_g41798 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_152, A2 => TL01_CLR1_n_164, ZN => TL01_CLR1_n_252);
  TL01_CLR1_g41799 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_163, A2 => char2perc(4), ZN => TL01_CLR1_n_251);
  TL01_CLR1_g41800 : NR2D0BWP7T port map(A1 => TL01_CLR1_n_164, A2 => char1perc(4), ZN => TL01_CLR1_n_250);
  TL01_CLR1_g41801 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_115, A2 => vcountintern(2), ZN => TL01_CLR1_n_249);
  TL01_CLR1_g41802 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_146, A2 => hcountintern(1), ZN => TL01_CLR1_n_248);
  TL01_CLR1_g41803 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_1495, A2 => hcountintern(1), ZN => TL01_CLR1_n_246);
  TL01_CLR1_g41804 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_185, A2 => TL01_CLR1_char2_sprite_frame_control_state_0, ZN => TL01_CLR1_n_1483);
  TL01_CLR1_g41805 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_139, A2 => FE_PHN106_TL01_CLR1_char1_sprite_frame_control_state_0, ZN => TL01_CLR1_n_1492);
  TL01_CLR1_g41806 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_162, A2 => char2perc(4), ZN => TL01_CLR1_n_242);
  TL01_CLR1_g41807 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_108, A2 => FE_DBTN12_char1perc_4, ZN => TL01_CLR1_n_240);
  TL01_CLR1_g41808 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_150, A2 => hcountintern(1), ZN => TL01_CLR1_n_238);
  TL01_CLR1_g41809 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_150, A2 => TL01_CLR1_n_85, ZN => TL01_CLR1_n_237);
  TL01_CLR1_g41810 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_103, A2 => hcountintern(1), ZN => TL01_CLR1_n_235);
  TL01_CLR1_g41811 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_145, A2 => hcountintern(1), ZN => TL01_CLR1_n_233);
  TL01_CLR1_g41812 : INVD0BWP7T port map(I => TL01_CLR1_n_222, ZN => TL01_CLR1_n_223);
  TL01_CLR1_g41813 : INVD0BWP7T port map(I => TL01_CLR1_n_219, ZN => TL01_CLR1_n_220);
  TL01_CLR1_g41814 : INVD0BWP7T port map(I => TL01_CLR1_n_208, ZN => TL01_CLR1_n_207);
  TL01_CLR1_g41815 : INVD0BWP7T port map(I => TL01_CLR1_n_206, ZN => TL01_CLR1_n_205);
  TL01_CLR1_g41816 : INVD0BWP7T port map(I => TL01_CLR1_n_200, ZN => TL01_CLR1_n_199);
  TL01_CLR1_g41817 : INVD1BWP7T port map(I => TL01_CLR1_n_198, ZN => TL01_CLR1_n_197);
  TL01_CLR1_g41818 : INVD1BWP7T port map(I => TL01_CLR1_n_194, ZN => TL01_CLR1_n_193);
  TL01_CLR1_g41819 : OAI21D0BWP7T port map(A1 => TL01_CLR1_char2_sprite_frame_control_frame_count_1, A2 => TL01_CLR1_char2_sprite_frame_control_frame_count_2, B => TL01_CLR1_char2_sprite_frame_control_frame_count_3, ZN => TL01_CLR1_n_189);
  TL01_CLR1_g41820 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_54, A2 => TL01_CLR1_n_90, B => hcountintern(8), ZN => TL01_CLR1_n_188);
  TL01_CLR1_g41821 : OR2D1BWP7T port map(A1 => TL01_CLR1_n_112, A2 => TL01_CLR1_n_77, Z => TL01_CLR1_n_187);
  TL01_CLR1_g41822 : OAI21D0BWP7T port map(A1 => TL01_CLR1_char1_sprite_frame_control_frame_count_1, A2 => FE_PHN111_TL01_CLR1_char1_sprite_frame_control_frame_count_2, B => FE_PHN109_TL01_CLR1_char1_sprite_frame_control_frame_count_3, ZN => TL01_CLR1_n_186);
  TL01_CLR1_g41823 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_121, B1 => TL01_CLR1_n_112, ZN => TL01_CLR1_n_227);
  TL01_CLR1_g41824 : INR2XD0BWP7T port map(A1 => TL01_CLR1_n_182, B1 => TL01_CLR1_n_129, ZN => TL01_CLR1_n_226);
  TL01_CLR1_g41825 : CKAN2D1BWP7T port map(A1 => TL01_CLR1_n_127, A2 => TL01_CLR1_n_136, Z => TL01_CLR1_n_225);
  TL01_CLR1_g41826 : NR3D0BWP7T port map(A1 => char2perc(4), A2 => char2perc(1), A3 => char2perc(0), ZN => TL01_CLR1_n_224);
  TL01_CLR1_g41827 : NR3D0BWP7T port map(A1 => char1perc(4), A2 => char1perc(1), A3 => char1perc(0), ZN => TL01_CLR1_n_222);
  TL01_CLR1_g41828 : AN2D0BWP7T port map(A1 => TL01_CLR1_n_138, A2 => char2perc(4), Z => TL01_CLR1_n_221);
  TL01_CLR1_g41829 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_146, A2 => TL01_CLR1_n_100, ZN => TL01_CLR1_n_219);
  TL01_CLR1_g41830 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_119, A2 => TL01_CLR1_n_111, ZN => TL01_CLR1_n_218);
  TL01_CLR1_g41831 : AOI21D0BWP7T port map(A1 => vcountintern(2), A2 => char1posy(1), B => TL01_CLR1_n_183, ZN => TL01_CLR1_n_217);
  TL01_CLR1_g41832 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_87, A2 => FE_DBTN13_char1perc_5, B1 => char1perc(6), B2 => char1perc(5), ZN => TL01_CLR1_n_216);
  TL01_CLR1_g41833 : OAI22D0BWP7T port map(A1 => vcountintern(2), A2 => char2posy(1), B1 => TL01_CLR1_n_57, B2 => TL01_CLR1_n_65, ZN => TL01_CLR1_n_215);
  TL01_CLR1_g41834 : NR4D0BWP7T port map(A1 => inputsp1(6), A2 => inputsp1(7), A3 => inputsp1(5), A4 => inputsp1(4), ZN => TL01_CLR1_n_214);
  TL01_CLR1_g41835 : NR4D0BWP7T port map(A1 => inputsp2(6), A2 => inputsp2(7), A3 => FE_PHN98_inputsp2_5, A4 => inputsp2(4), ZN => TL01_CLR1_n_213);
  TL01_CLR1_g41836 : MOAI22D0BWP7T port map(A1 => FE_DBTN1_char2posx_1, A2 => char2posx(2), B1 => FE_DBTN1_char2posx_1, B2 => char2posx(2), ZN => TL01_CLR1_n_212);
  TL01_CLR1_g41837 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_66, A2 => char1posx(2), B1 => TL01_CLR1_n_66, B2 => char1posx(2), ZN => TL01_CLR1_n_211);
  TL01_CLR1_g41839 : AOI22D0BWP7T port map(A1 => TL01_CLR1_n_92, A2 => vcountintern(2), B1 => TL01_CLR1_n_57, B2 => vcountintern(1), ZN => TL01_CLR1_n_209);
  TL01_CLR1_g41840 : XNR2D1BWP7T port map(A1 => inputsp1(1), A2 => inputsp1(0), ZN => TL01_CLR1_n_208);
  TL01_CLR1_g41841 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_154, A2 => hcountintern(9), ZN => TL01_CLR1_n_206);
  TL01_CLR1_g41842 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_65, A2 => char2posy(2), B1 => TL01_CLR1_n_65, B2 => char2posy(2), ZN => TL01_CLR1_n_204);
  TL01_CLR1_g41843 : AOI21D0BWP7T port map(A1 => char2posy(0), A2 => char2posy(1), B => char2posy(2), ZN => TL01_CLR1_n_203);
  TL01_CLR1_g41844 : CKXOR2D1BWP7T port map(A1 => inputsp2(1), A2 => inputsp2(0), Z => TL01_CLR1_n_202);
  TL01_CLR1_g41845 : AOI21D0BWP7T port map(A1 => FE_DBTN10_char1perc_1, A2 => char1perc(5), B => TL01_CLR1_n_133, ZN => TL01_CLR1_n_201);
  TL01_CLR1_g41846 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_105, A2 => TL01_CLR1_n_113, ZN => TL01_CLR1_n_200);
  TL01_CLR1_g41847 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_103, A2 => TL01_CLR1_n_113, ZN => TL01_CLR1_n_198);
  TL01_CLR1_g41848 : AOI21D0BWP7T port map(A1 => FE_DBTN5_char2perc_1, A2 => char2perc(5), B => TL01_CLR1_n_134, ZN => TL01_CLR1_n_196);
  TL01_CLR1_g41849 : AOI21D0BWP7T port map(A1 => char1posy(0), A2 => char1posy(1), B => char1posy(2), ZN => TL01_CLR1_n_195);
  TL01_CLR1_g41850 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_104, A2 => TL01_CLR1_n_149, ZN => TL01_CLR1_n_194);
  TL01_CLR1_g41851 : OAI22D0BWP7T port map(A1 => TL01_CLR1_n_77, A2 => char2perc(3), B1 => FE_DBTN7_char2perc_3, B2 => char2perc(7), ZN => TL01_CLR1_n_192);
  TL01_CLR1_g41852 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_56, A2 => char1perc(3), B => TL01_CLR1_n_178, ZN => TL01_CLR1_n_191);
  TL01_CLR1_g41853 : AOI21D0BWP7T port map(A1 => TL01_CLR1_n_55, A2 => vcountintern(1), B => TL01_CLR1_n_116, ZN => TL01_CLR1_n_190);
  TL01_CLR1_g41854 : INVD1BWP7T port map(I => TL01_CLR1_n_171, ZN => TL01_CLR1_n_170);
  TL01_CLR1_g41855 : INVD0BWP7T port map(I => TL01_CLR1_n_168, ZN => TL01_CLR1_n_167);
  TL01_CLR1_g41856 : INVD0BWP7T port map(I => TL01_CLR1_n_166, ZN => TL01_CLR1_n_165);
  TL01_CLR1_g41857 : INVD1BWP7T port map(I => TL01_CLR1_n_162, ZN => TL01_CLR1_n_161);
  TL01_CLR1_g41858 : INVD1BWP7T port map(I => TL01_CLR1_n_160, ZN => TL01_CLR1_n_1494);
  TL01_CLR1_g41859 : INVD0BWP7T port map(I => TL01_CLR1_n_158, ZN => TL01_CLR1_n_157);
  TL01_CLR1_g41860 : INVD1BWP7T port map(I => TL01_CLR1_n_156, ZN => TL01_CLR1_n_155);
  TL01_CLR1_g41861 : INVD0BWP7T port map(I => TL01_CLR1_n_154, ZN => TL01_CLR1_n_153);
  TL01_CLR1_g41862 : INVD1BWP7T port map(I => TL01_CLR1_n_152, ZN => TL01_CLR1_n_151);
  TL01_CLR1_g41863 : INVD0BWP7T port map(I => TL01_CLR1_n_150, ZN => TL01_CLR1_n_149);
  TL01_CLR1_g41864 : INVD1BWP7T port map(I => TL01_CLR1_n_148, ZN => TL01_CLR1_n_147);
  TL01_CLR1_g41865 : INVD1BWP7T port map(I => TL01_CLR1_n_146, ZN => TL01_CLR1_n_145);
  TL01_CLR1_g41866 : NR2XD0BWP7T port map(A1 => char2posy(0), A2 => char2posy(1), ZN => TL01_CLR1_n_144);
  TL01_CLR1_g41867 : INR2D1BWP7T port map(A1 => TL01_CLR1_char2_sprite_frame_control_state_1, B1 => FE_PHN99_TL01_CLR1_char2_sprite_frame_control_state_2, ZN => TL01_CLR1_n_185);
  TL01_CLR1_g41868 : NR2XD0BWP7T port map(A1 => vcountintern(1), A2 => vcountintern(2), ZN => TL01_CLR1_n_184);
  TL01_CLR1_g41869 : NR2XD0BWP7T port map(A1 => vcountintern(2), A2 => char1posy(1), ZN => TL01_CLR1_n_183);
  TL01_CLR1_g41870 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_87, A2 => char1perc(2), ZN => TL01_CLR1_n_182);
  TL01_CLR1_g41871 : OR2D1BWP7T port map(A1 => TL01_CLR1_char1_sprite_frame_control_state_0, A2 => TL01_CLR1_char1_sprite_frame_control_state_1, Z => TL01_CLR1_n_1491);
  TL01_CLR1_g41872 : ND2D1BWP7T port map(A1 => TL01_CLR1_char1_sprite_frame_control_frame_count_1, A2 => TL01_CLR1_char1_sprite_frame_control_frame_count_0, ZN => TL01_CLR1_n_1487);
  TL01_CLR1_g41873 : ND2D1BWP7T port map(A1 => char2posx(0), A2 => char2posx(1), ZN => TL01_CLR1_n_181);
  TL01_CLR1_g41874 : ND2D1BWP7T port map(A1 => TL01_CLR1_char2_sprite_frame_control_frame_count_1, A2 => TL01_CLR1_char2_sprite_frame_control_frame_count_0, ZN => TL01_CLR1_n_1478);
  TL01_CLR1_g41875 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_85, A2 => char2posx(0), ZN => TL01_CLR1_n_143);
  TL01_CLR1_g41876 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_85, A2 => char1posx(0), ZN => TL01_CLR1_n_142);
  TL01_CLR1_g41877 : OR2D1BWP7T port map(A1 => TL01_CLR1_char1_sprite_frame_control_state_2, A2 => TL01_CLR1_char1_sprite_frame_control_state_1, Z => TL01_CLR1_n_1490);
  TL01_CLR1_g41878 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_92, A2 => char2posy(0), ZN => TL01_CLR1_n_180);
  TL01_CLR1_g41879 : NR2D1BWP7T port map(A1 => FE_DBTN13_char1perc_5, A2 => char1perc(3), ZN => TL01_CLR1_n_179);
  TL01_CLR1_g41880 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_56, A2 => char1perc(3), ZN => TL01_CLR1_n_178);
  TL01_CLR1_g41881 : ND2D1BWP7T port map(A1 => char1posx(1), A2 => char1posx(2), ZN => TL01_CLR1_n_177);
  TL01_CLR1_g41882 : NR2XD0BWP7T port map(A1 => vcountintern(4), A2 => vcountintern(5), ZN => TL01_CLR1_n_176);
  TL01_CLR1_g41883 : NR2D0BWP7T port map(A1 => char1perc(5), A2 => char1perc(1), ZN => TL01_CLR1_n_175);
  TL01_CLR1_g41884 : NR2D0BWP7T port map(A1 => char2perc(5), A2 => char2perc(1), ZN => TL01_CLR1_n_174);
  TL01_CLR1_g41885 : NR2XD0BWP7T port map(A1 => char2perc(4), A2 => char2perc(3), ZN => TL01_CLR1_n_173);
  TL01_CLR1_g41886 : ND2D1BWP7T port map(A1 => char2perc(5), A2 => char2perc(1), ZN => TL01_CLR1_n_172);
  TL01_CLR1_g41887 : ND2D1BWP7T port map(A1 => char1perc(5), A2 => char1perc(1), ZN => TL01_CLR1_n_171);
  TL01_CLR1_g41888 : AN2D1BWP7T port map(A1 => vcountintern(7), A2 => vcountintern(6), Z => TL01_CLR1_n_169);
  TL01_CLR1_g41889 : CKND2D1BWP7T port map(A1 => TL01_CLR1_n_53, A2 => TL01_CLR1_n_84, ZN => TL01_CLR1_n_168);
  TL01_CLR1_g41890 : NR2D1BWP7T port map(A1 => hcountintern(8), A2 => hcountintern(9), ZN => TL01_CLR1_n_166);
  TL01_CLR1_g41891 : CKND2D1BWP7T port map(A1 => char1perc(6), A2 => char1perc(2), ZN => TL01_CLR1_n_164);
  TL01_CLR1_g41892 : CKND2D1BWP7T port map(A1 => char2perc(6), A2 => char2perc(2), ZN => TL01_CLR1_n_163);
  TL01_CLR1_g41893 : NR2D1BWP7T port map(A1 => char2perc(6), A2 => char2perc(2), ZN => TL01_CLR1_n_162);
  TL01_CLR1_g41894 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_83, A2 => TL01_CLR1_n_86, ZN => TL01_CLR1_n_160);
  TL01_CLR1_g41895 : ND2D1BWP7T port map(A1 => vcountintern(1), A2 => vcountintern(2), ZN => TL01_CLR1_n_159);
  TL01_CLR1_g41896 : ND2D1BWP7T port map(A1 => hcountintern(6), A2 => hcountintern(7), ZN => TL01_CLR1_n_158);
  TL01_CLR1_g41897 : CKND2D1BWP7T port map(A1 => TL01_CLR1_n_56, A2 => FE_DBTN11_char1perc_3, ZN => TL01_CLR1_n_156);
  TL01_CLR1_g41898 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_90, A2 => TL01_CLR1_n_82, ZN => TL01_CLR1_n_154);
  TL01_CLR1_g41899 : ND2D1BWP7T port map(A1 => char1perc(7), A2 => char1perc(3), ZN => TL01_CLR1_n_152);
  TL01_CLR1_g41900 : NR2XD0BWP7T port map(A1 => hcountintern(3), A2 => hcountintern(2), ZN => TL01_CLR1_n_150);
  TL01_CLR1_g41901 : NR2D1BWP7T port map(A1 => vcountintern(8), A2 => vcountintern(9), ZN => TL01_CLR1_n_148);
  TL01_CLR1_g41902 : CKND2D1BWP7T port map(A1 => hcountintern(3), A2 => hcountintern(2), ZN => TL01_CLR1_n_146);
  TL01_CLR1_g41903 : INVD0BWP7T port map(I => TL01_CLR1_n_135, ZN => TL01_CLR1_n_1482);
  TL01_CLR1_g41904 : INVD0BWP7T port map(I => TL01_CLR1_n_1563, ZN => TL01_CLR1_n_123);
  TL01_CLR1_g41905 : INVD0BWP7T port map(I => TL01_CLR1_n_117, ZN => TL01_CLR1_n_1481);
  TL01_CLR1_g41906 : INVD0BWP7T port map(I => TL01_CLR1_n_115, ZN => TL01_CLR1_n_114);
  TL01_CLR1_g41907 : INVD1BWP7T port map(I => TL01_CLR1_n_111, ZN => TL01_CLR1_n_110);
  TL01_CLR1_g41908 : INVD1BWP7T port map(I => TL01_CLR1_n_109, ZN => TL01_CLR1_n_108);
  TL01_CLR1_g41909 : INVD1BWP7T port map(I => TL01_CLR1_n_107, ZN => TL01_CLR1_n_106);
  TL01_CLR1_g41910 : INVD1BWP7T port map(I => TL01_CLR1_n_105, ZN => TL01_CLR1_n_104);
  TL01_CLR1_g41911 : INVD1BWP7T port map(I => TL01_CLR1_n_1495, ZN => TL01_CLR1_n_103);
  TL01_CLR1_g41912 : INVD1BWP7T port map(I => TL01_CLR1_n_101, ZN => TL01_CLR1_n_100);
  TL01_CLR1_g41913 : INR2D1BWP7T port map(A1 => char1posy(0), B1 => vcountintern(1), ZN => TL01_CLR1_n_141);
  TL01_CLR1_g41914 : CKND2D1BWP7T port map(A1 => FE_DBTN8_char2perc_4, A2 => char2perc(5), ZN => TL01_CLR1_n_140);
  TL01_CLR1_g41915 : INR2D1BWP7T port map(A1 => TL01_CLR1_char1_sprite_frame_control_state_1, B1 => TL01_CLR1_char1_sprite_frame_control_state_2, ZN => TL01_CLR1_n_139);
  TL01_CLR1_g41916 : CKND2D1BWP7T port map(A1 => FE_DBTN7_char2perc_3, A2 => char2perc(5), ZN => TL01_CLR1_n_138);
  TL01_CLR1_g41917 : CKND2D1BWP7T port map(A1 => char1posx(1), A2 => char1posx(0), ZN => TL01_CLR1_n_137);
  TL01_CLR1_g41918 : CKND2D1BWP7T port map(A1 => TL01_CLR1_n_61, A2 => char2perc(2), ZN => TL01_CLR1_n_136);
  TL01_CLR1_g41919 : NR2D1BWP7T port map(A1 => TL01_CLR1_char2_sprite_frame_control_state_0, A2 => TL01_CLR1_char2_sprite_frame_control_state_1, ZN => TL01_CLR1_n_135);
  TL01_CLR1_g41920 : NR2D1BWP7T port map(A1 => FE_DBTN5_char2perc_1, A2 => char2perc(5), ZN => TL01_CLR1_n_134);
  TL01_CLR1_g41921 : NR2D1BWP7T port map(A1 => FE_DBTN10_char1perc_1, A2 => char1perc(5), ZN => TL01_CLR1_n_133);
  TL01_CLR1_g41922 : NR2D1BWP7T port map(A1 => char1perc(4), A2 => char1perc(3), ZN => TL01_CLR1_n_132);
  TL01_CLR1_g41923 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_56, A2 => char1perc(6), ZN => TL01_CLR1_n_131);
  TL01_CLR1_g41924 : NR2D0BWP7T port map(A1 => char1perc(6), A2 => char1perc(4), ZN => TL01_CLR1_n_130);
  TL01_CLR1_g41925 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_87, A2 => char1perc(2), ZN => TL01_CLR1_n_129);
  TL01_CLR1_g41926 : CKAN2D1BWP7T port map(A1 => char2posy(1), A2 => char2posy(2), Z => TL01_CLR1_n_128);
  TL01_CLR1_g41927 : CKND2D1BWP7T port map(A1 => FE_DBTN6_char2perc_2, A2 => char2perc(6), ZN => TL01_CLR1_n_127);
  TL01_CLR1_g41928 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_52, A2 => vcountintern(0), ZN => TL01_CLR1_n_126);
  TL01_CLR1_g41929 : CKND2D1BWP7T port map(A1 => char1posy(2), A2 => char1posy(1), ZN => TL01_CLR1_n_125);
  TL01_CLR1_g41930 : NR2D1BWP7T port map(A1 => hcountintern(4), A2 => TL01_CLR1_n_84, ZN => TL01_CLR1_n_124);
  TL01_CLR1_g41932 : ND2D1BWP7T port map(A1 => hcountintern(4), A2 => TL01_CLR1_n_84, ZN => TL01_CLR1_n_1493);
  TL01_CLR1_g41933 : CKND2D1BWP7T port map(A1 => TL01_CLR1_n_77, A2 => char2perc(6), ZN => TL01_CLR1_n_121);
  TL01_CLR1_g41934 : NR2D1BWP7T port map(A1 => FE_DBTN9_char2perc_5, A2 => char2perc(6), ZN => TL01_CLR1_n_120);
  TL01_CLR1_g41935 : ND2D1BWP7T port map(A1 => TL01_CLR1_n_56, A2 => char1perc(6), ZN => TL01_CLR1_n_119);
  TL01_CLR1_g41936 : CKND2D1BWP7T port map(A1 => char2posx(2), A2 => char2posx(1), ZN => TL01_CLR1_n_118);
  TL01_CLR1_g41937 : NR2D1BWP7T port map(A1 => FE_PHN99_TL01_CLR1_char2_sprite_frame_control_state_2, A2 => TL01_CLR1_char2_sprite_frame_control_state_1, ZN => TL01_CLR1_n_117);
  TL01_CLR1_g41938 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_55, A2 => vcountintern(1), ZN => TL01_CLR1_n_116);
  TL01_CLR1_g41939 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_55, A2 => TL01_CLR1_n_92, ZN => TL01_CLR1_n_115);
  TL01_CLR1_g41940 : NR2XD0BWP7T port map(A1 => hcountintern(1), A2 => TL01_hcount_int(0), ZN => TL01_CLR1_n_113);
  TL01_CLR1_g41941 : NR2D1BWP7T port map(A1 => char2perc(4), A2 => char2perc(5), ZN => TL01_CLR1_n_112);
  TL01_CLR1_g41942 : ND2D1BWP7T port map(A1 => FE_DBTN13_char1perc_5, A2 => FE_DBTN12_char1perc_4, ZN => TL01_CLR1_n_111);
  TL01_CLR1_g41943 : NR2D1BWP7T port map(A1 => char1perc(6), A2 => char1perc(2), ZN => TL01_CLR1_n_109);
  TL01_CLR1_g41944 : NR2XD0BWP7T port map(A1 => vcountintern(6), A2 => vcountintern(7), ZN => TL01_CLR1_n_107);
  TL01_CLR1_g41945 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_85, A2 => TL01_CLR1_n_51, ZN => TL01_CLR1_n_105);
  TL01_CLR1_g41946 : CKND2D1BWP7T port map(A1 => TL01_CLR1_n_54, A2 => hcountintern(2), ZN => TL01_CLR1_n_1495);
  TL01_CLR1_g41947 : ND2D1BWP7T port map(A1 => FE_DBTN7_char2perc_3, A2 => TL01_CLR1_n_77, ZN => TL01_CLR1_n_102);
  TL01_CLR1_g41948 : NR2XD0BWP7T port map(A1 => TL01_CLR1_n_84, A2 => TL01_CLR1_n_53, ZN => TL01_CLR1_n_101);
  TL01_CLR1_g41949 : CKND2D1BWP7T port map(A1 => char2perc(3), A2 => char2perc(7), ZN => TL01_CLR1_n_99);
  TL01_CLR1_g41950 : INVD1BWP7T port map(I => char2posy(6), ZN => TL01_CLR1_n_98);
  TL01_CLR1_g41951 : INVD0BWP7T port map(I => inputsp1(3), ZN => TL01_CLR1_n_97);
  TL01_CLR1_g41953 : INVD0BWP7T port map(I => inputsp1(2), ZN => TL01_CLR1_n_95);
  TL01_CLR1_g41956 : INVD0BWP7T port map(I => vcountintern(1), ZN => TL01_CLR1_n_92);
  TL01_CLR1_g41958 : INVD0BWP7T port map(I => hcountintern(6), ZN => TL01_CLR1_n_90);
  TL01_CLR1_g41961 : INVD1BWP7T port map(I => char1perc(6), ZN => TL01_CLR1_n_87);
  TL01_CLR1_g41962 : INVD1BWP7T port map(I => vcountintern(5), ZN => TL01_CLR1_n_86);
  TL01_CLR1_g41963 : INVD1BWP7T port map(I => hcountintern(1), ZN => TL01_CLR1_n_85);
  TL01_CLR1_g41964 : INVD1BWP7T port map(I => hcountintern(5), ZN => TL01_CLR1_n_84);
  TL01_CLR1_g41965 : INVD1BWP7T port map(I => vcountintern(4), ZN => TL01_CLR1_n_83);
  TL01_CLR1_g41966 : INVD1BWP7T port map(I => hcountintern(7), ZN => TL01_CLR1_n_82);
  TL01_CLR1_g41967 : INVD1BWP7T port map(I => hcountintern(9), ZN => TL01_CLR1_n_81);
  TL01_CLR1_g41971 : INVD1BWP7T port map(I => char2perc(7), ZN => TL01_CLR1_n_77);
  TL01_CLR1_g41973 : INVD0BWP7T port map(I => char2posx(4), ZN => TL01_CLR1_n_75);
  TL01_CLR1_g41974 : INVD1BWP7T port map(I => char1posy(6), ZN => TL01_CLR1_n_74);
  TL01_CLR1_g41975 : CKND1BWP7T port map(I => inputsp2(2), ZN => TL01_CLR1_n_73);
  TL01_CLR1_g41976 : INVD0BWP7T port map(I => orientationp1, ZN => TL01_CLR1_n_72);
  TL01_CLR1_g41977 : INVD1BWP7T port map(I => orientationp2, ZN => TL01_CLR1_n_71);
  TL01_CLR1_g41979 : INVD0BWP7T port map(I => char1posx(0), ZN => TL01_CLR1_n_69);
  TL01_CLR1_g41980 : INVD0BWP7T port map(I => vcountintern(9), ZN => TL01_CLR1_n_68);
  TL01_CLR1_g41982 : INVD0BWP7T port map(I => char1posx(1), ZN => TL01_CLR1_n_66);
  TL01_CLR1_g41983 : INVD0BWP7T port map(I => char2posy(1), ZN => TL01_CLR1_n_65);
  TL01_CLR1_g41987 : INVD1BWP7T port map(I => char2perc(6), ZN => TL01_CLR1_n_61);
  TL01_CLR1_g41988 : INVD0BWP7T port map(I => hcountintern(8), ZN => TL01_CLR1_n_60);
  TL01_CLR1_g41989 : INVD1BWP7T port map(I => vcountintern(7), ZN => TL01_CLR1_n_59);
  TL01_CLR1_g41991 : INVD1BWP7T port map(I => vcountintern(2), ZN => TL01_CLR1_n_57);
  TL01_CLR1_g41992 : INVD1BWP7T port map(I => char1perc(7), ZN => TL01_CLR1_n_56);
  TL01_CLR1_g41993 : INVD1BWP7T port map(I => vcountintern(0), ZN => TL01_CLR1_n_55);
  TL01_CLR1_g41994 : INVD1BWP7T port map(I => hcountintern(3), ZN => TL01_CLR1_n_54);
  TL01_CLR1_g41995 : INVD1BWP7T port map(I => hcountintern(4), ZN => TL01_CLR1_n_53);
  TL01_CLR1_g41996 : INVD1BWP7T port map(I => vcountintern(3), ZN => TL01_CLR1_n_52);
  TL01_CLR1_g41997 : INVD1BWP7T port map(I => TL01_hcount_int(0), ZN => TL01_CLR1_n_51);
  TL01_CLR1_char1_sprite_frame_control_sprite_reg_0 : DFKCND1BWP7T port map(CN => FE_DBTN14_reset, CP => CTS_16, D => TL01_CLR1_n_305, Q => TL01_CLR1_char1_sprite_sprite_0, QN => TL01_CLR1_n_50);
  TL01_CLR1_g2 : IIND4D0BWP7T port map(A1 => TL01_CLR1_n_1418, A2 => TL01_CLR1_n_1429, B1 => TL01_CLR1_n_1445, B2 => TL01_CLR1_n_1426, ZN => TL01_CLR1_n_49);
  TL01_CLR1_g42000 : INR2D1BWP7T port map(A1 => TL01_CLR1_n_1110, B1 => TL01_CLR1_n_800, ZN => TL01_CLR1_n_48);
  TL01_CLR1_g42001 : IINR4D0BWP7T port map(A1 => TL01_CLR1_n_1341, A2 => TL01_CLR1_n_1017, B1 => TL01_CLR1_n_1226, B2 => TL01_CLR1_n_1277, ZN => TL01_CLR1_n_47);
  TL01_CLR1_g42002 : INR3D0BWP7T port map(A1 => TL01_CLR1_n_967, B1 => TL01_CLR1_n_731, B2 => TL01_CLR1_n_757, ZN => TL01_CLR1_n_46);
  TL01_CLR1_g42003 : INR3D0BWP7T port map(A1 => TL01_CLR1_n_729, B1 => TL01_CLR1_n_975, B2 => TL01_CLR1_n_959, ZN => TL01_CLR1_n_45);
  TL01_CLR1_g42004 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_643, B1 => vcountintern(0), ZN => TL01_CLR1_n_44);
  TL01_CLR1_g42005 : INR2D1BWP7T port map(A1 => TL01_CLR1_n_283, B1 => TL01_CLR1_n_600, ZN => TL01_CLR1_n_43);
  TL01_CLR1_g42006 : IIND4D0BWP7T port map(A1 => TL01_CLR1_n_264, A2 => TL01_CLR1_n_267, B1 => TL01_CLR1_n_428, B2 => TL01_CLR1_n_435, ZN => TL01_CLR1_n_42);
  TL01_CLR1_char1_sprite_frame_control_cnt_cur_count_reg_4 : DFKCNQD1BWP7T port map(CN => FE_PHN59_TL01_CLR1_char1_sprite_frame_control_cnt_reset, CP => CTS_16, D => TL01_CLR1_n_40, Q => FE_PHN105_TL01_CLR1_char1_sprite_frame_control_frame_count_4);
  TL01_CLR1_char2_sprite_frame_control_cnt_cur_count_reg_4 : DFKCNQD1BWP7T port map(CN => FE_PHN169_TL01_CLR1_char2_sprite_frame_control_cnt_reset, CP => CTS_15, D => FE_PHN153_TL01_CLR1_n_41, Q => TL01_CLR1_char2_sprite_frame_control_frame_count_4);
  TL01_CLR1_char2_sprite_frame_control_cnt_cur_count_reg_3 : DFKCNQD1BWP7T port map(CN => FE_PHN169_TL01_CLR1_char2_sprite_frame_control_cnt_reset, CP => CTS_15, D => TL01_CLR1_n_39, Q => TL01_CLR1_char2_sprite_frame_control_frame_count_3);
  TL01_CLR1_char1_sprite_frame_control_cnt_cur_count_reg_3 : DFKCNQD1BWP7T port map(CN => FE_PHN59_TL01_CLR1_char1_sprite_frame_control_cnt_reset, CP => CTS_16, D => TL01_CLR1_n_37, Q => TL01_CLR1_char1_sprite_frame_control_frame_count_3);
  TL01_CLR1_g1919 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_29, A2 => TL01_CLR1_n_38, B1 => TL01_CLR1_n_29, B2 => FE_PHN163_TL01_CLR1_char2_sprite_frame_control_frame_count_4, ZN => TL01_CLR1_n_41);
  TL01_CLR1_g1920 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_29, A2 => TL01_CLR1_n_36, B1 => TL01_CLR1_n_29, B2 => TL01_CLR1_char1_sprite_frame_control_frame_count_4, ZN => TL01_CLR1_n_40);
  TL01_CLR1_char2_sprite_frame_control_cnt_cur_count_reg_1 : DFKCNQD1BWP7T port map(CN => FE_PHN169_TL01_CLR1_char2_sprite_frame_control_cnt_reset, CP => CTS_15, D => FE_PHN150_TL01_CLR1_n_34, Q => TL01_CLR1_char2_sprite_frame_control_frame_count_1);
  TL01_CLR1_char1_sprite_frame_control_cnt_cur_count_reg_1 : DFKCNQD1BWP7T port map(CN => FE_PHN59_TL01_CLR1_char1_sprite_frame_control_cnt_reset, CP => CTS_16, D => TL01_CLR1_n_32, Q => TL01_CLR1_char1_sprite_frame_control_frame_count_1);
  TL01_CLR1_char2_sprite_frame_control_cnt_cur_count_reg_2 : DFKCNQD1BWP7T port map(CN => FE_PHN169_TL01_CLR1_char2_sprite_frame_control_cnt_reset, CP => CTS_15, D => FE_PHN154_TL01_CLR1_n_33, Q => TL01_CLR1_char2_sprite_frame_control_frame_count_2);
  TL01_CLR1_char1_sprite_frame_control_cnt_cur_count_reg_2 : DFKCNQD1BWP7T port map(CN => FE_PHN59_TL01_CLR1_char1_sprite_frame_control_cnt_reset, CP => CTS_16, D => TL01_CLR1_n_31, Q => TL01_CLR1_char1_sprite_frame_control_frame_count_2);
  TL01_CLR1_char1_sprite_frame_control_cnt_cur_count_reg_0 : DFKCNQD1BWP7T port map(CN => FE_PHN59_TL01_CLR1_char1_sprite_frame_control_cnt_reset, CP => CTS_16, D => TL01_CLR1_n_30, Q => FE_PHN108_TL01_CLR1_char1_sprite_frame_control_frame_count_0);
  TL01_CLR1_char2_sprite_frame_control_cnt_cur_count_reg_0 : DFKCNQD1BWP7T port map(CN => FE_PHN169_TL01_CLR1_char2_sprite_frame_control_cnt_reset, CP => CTS_15, D => TL01_CLR1_n_35, Q => FE_PHN107_TL01_CLR1_char2_sprite_frame_control_frame_count_0);
  TL01_CLR1_g1927 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_29, A2 => TL01_CLR1_n_26, B1 => TL01_CLR1_n_29, B2 => FE_PHN84_TL01_CLR1_char2_sprite_frame_control_frame_count_3, ZN => TL01_CLR1_n_39);
  TL01_CLR1_char2_sprite_frame_control_cnt_reset_reg : DFXD1BWP7T port map(CP => CTS_15, DA => FE_PHN53_TL01_CLR1_n_1, DB => TL01_CLR1_n_28, Q => TL01_CLR1_n_1, QN => TL01_CLR1_char2_sprite_frame_control_cnt_reset, SA => FE_OFN3_reset);
  TL01_CLR1_char1_sprite_frame_control_cnt_reset_reg : DFXD1BWP7T port map(CP => CTS_16, DA => TL01_CLR1_n_0, DB => TL01_CLR1_n_27, Q => FE_PHN51_TL01_CLR1_n_0, QN => TL01_CLR1_char1_sprite_frame_control_cnt_reset, SA => FE_OFN3_reset);
  TL01_CLR1_g1930 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_24, A2 => TL01_CLR1_char2_sprite_frame_control_frame_count_4, B1 => TL01_CLR1_n_24, B2 => TL01_CLR1_char2_sprite_frame_control_frame_count_4, ZN => TL01_CLR1_n_38);
  TL01_CLR1_g1931 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_29, A2 => TL01_CLR1_n_25, B1 => TL01_CLR1_n_29, B2 => FE_PHN109_TL01_CLR1_char1_sprite_frame_control_frame_count_3, ZN => TL01_CLR1_n_37);
  TL01_CLR1_g1932 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_23, A2 => TL01_CLR1_char1_sprite_frame_control_frame_count_4, B1 => TL01_CLR1_n_23, B2 => TL01_CLR1_char1_sprite_frame_control_frame_count_4, ZN => TL01_CLR1_n_36);
  TL01_CLR1_g1933 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_29, A2 => TL01_CLR1_char2_sprite_frame_control_frame_count_0, B1 => TL01_CLR1_n_29, B2 => TL01_CLR1_char2_sprite_frame_control_frame_count_0, ZN => TL01_CLR1_n_35);
  TL01_CLR1_g1934 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_29, A2 => TL01_CLR1_n_14, B1 => TL01_CLR1_n_29, B2 => TL01_CLR1_char2_sprite_frame_control_frame_count_1, ZN => TL01_CLR1_n_34);
  TL01_CLR1_g1935 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_29, A2 => TL01_CLR1_n_15, B1 => TL01_CLR1_n_29, B2 => FE_PHN171_TL01_CLR1_char2_sprite_frame_control_frame_count_2, ZN => TL01_CLR1_n_33);
  TL01_CLR1_g1936 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_29, A2 => TL01_CLR1_n_12, B1 => TL01_CLR1_n_29, B2 => TL01_CLR1_char1_sprite_frame_control_frame_count_1, ZN => FE_PHN151_TL01_CLR1_n_32);
  TL01_CLR1_g1937 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_29, A2 => TL01_CLR1_n_11, B1 => TL01_CLR1_n_29, B2 => FE_PHN111_TL01_CLR1_char1_sprite_frame_control_frame_count_2, ZN => TL01_CLR1_n_31);
  TL01_CLR1_g1938 : MOAI22D0BWP7T port map(A1 => TL01_CLR1_n_29, A2 => FE_PHN161_TL01_CLR1_char1_sprite_frame_control_frame_count_0, B1 => TL01_CLR1_n_29, B2 => TL01_CLR1_char1_sprite_frame_control_frame_count_0, ZN => TL01_CLR1_n_30);
  TL01_CLR1_g1939 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_1481, A2 => TL01_CLR1_n_1564, B => TL01_CLR1_n_17, C => TL01_CLR1_n_22, ZN => TL01_CLR1_n_28);
  TL01_CLR1_g1940 : IND4D1BWP7T port map(A1 => TL01_CLR1_n_13, B1 => TL01_CLR1_n_19, B2 => TL01_CLR1_n_16, B3 => TL01_CLR1_n_20, ZN => TL01_CLR1_n_29);
  TL01_CLR1_g1941 : OAI211D1BWP7T port map(A1 => TL01_CLR1_n_1490, A2 => TL01_CLR1_n_1565, B => TL01_CLR1_n_18, C => TL01_CLR1_n_21, ZN => TL01_CLR1_n_27);
  TL01_CLR1_g1942 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_9, A2 => FE_PHN84_TL01_CLR1_char2_sprite_frame_control_frame_count_3, B1 => TL01_CLR1_n_9, B2 => FE_PHN84_TL01_CLR1_char2_sprite_frame_control_frame_count_3, ZN => TL01_CLR1_n_26);
  TL01_CLR1_g1943 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_10, A2 => FE_PHN109_TL01_CLR1_char1_sprite_frame_control_frame_count_3, B1 => TL01_CLR1_n_10, B2 => FE_PHN109_TL01_CLR1_char1_sprite_frame_control_frame_count_3, ZN => TL01_CLR1_n_25);
  TL01_CLR1_g1944 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_9, B1 => FE_PHN84_TL01_CLR1_char2_sprite_frame_control_frame_count_3, ZN => TL01_CLR1_n_24);
  TL01_CLR1_g1945 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_10, B1 => FE_PHN109_TL01_CLR1_char1_sprite_frame_control_frame_count_3, ZN => TL01_CLR1_n_23);
  TL01_CLR1_g1946 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_5, A2 => FE_PHN99_TL01_CLR1_char2_sprite_frame_control_state_2, B => TL01_CLR1_n_1482, ZN => TL01_CLR1_n_22);
  TL01_CLR1_g1947 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_6, A2 => TL01_CLR1_char1_sprite_frame_control_state_2, B => FE_PHN172_TL01_CLR1_n_1491, ZN => TL01_CLR1_n_21);
  TL01_CLR1_g1948 : NR4D0BWP7T port map(A1 => TL01_CLR1_n_1493, A2 => TL01_CLR1_n_1494, A3 => TL01_CLR1_n_1495, A4 => TL01_CLR1_n_1563, ZN => TL01_CLR1_n_20);
  TL01_CLR1_g1949 : INR4D0BWP7T port map(A1 => hcountintern(1), B1 => TL01_hcount_int(0), B2 => hcountintern(7), B3 => hcountintern(6), ZN => TL01_CLR1_n_19);
  TL01_CLR1_g1950 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_3, A2 => TL01_CLR1_char1_sprite_frame_control_state_2, B => TL01_CLR1_n_1484, ZN => TL01_CLR1_n_18);
  TL01_CLR1_g1951 : OAI21D0BWP7T port map(A1 => TL01_CLR1_n_2, A2 => FE_PHN99_TL01_CLR1_char2_sprite_frame_control_state_2, B => TL01_CLR1_n_1475, ZN => TL01_CLR1_n_17);
  TL01_CLR1_g1952 : INR4D0BWP7T port map(A1 => vcountintern(2), B1 => vcountintern(1), B2 => vcountintern(0), B3 => vcountintern(3), ZN => TL01_CLR1_n_16);
  TL01_CLR1_g1953 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_1478, A2 => TL01_CLR1_char2_sprite_frame_control_frame_count_2, B1 => TL01_CLR1_n_1478, B2 => TL01_CLR1_char2_sprite_frame_control_frame_count_2, ZN => TL01_CLR1_n_15);
  TL01_CLR1_g1954 : XNR2D1BWP7T port map(A1 => TL01_CLR1_char2_sprite_frame_control_frame_count_0, A2 => TL01_CLR1_char2_sprite_frame_control_frame_count_1, ZN => TL01_CLR1_n_14);
  TL01_CLR1_g1955 : IND4D0BWP7T port map(A1 => vcountintern(9), B1 => vcountintern(8), B2 => vcountintern(6), B3 => vcountintern(7), ZN => TL01_CLR1_n_13);
  TL01_CLR1_g1956 : XNR2D1BWP7T port map(A1 => TL01_CLR1_char1_sprite_frame_control_frame_count_0, A2 => TL01_CLR1_char1_sprite_frame_control_frame_count_1, ZN => TL01_CLR1_n_12);
  TL01_CLR1_g1957 : MAOI22D0BWP7T port map(A1 => TL01_CLR1_n_1487, A2 => FE_PHN111_TL01_CLR1_char1_sprite_frame_control_frame_count_2, B1 => TL01_CLR1_n_1487, B2 => FE_PHN111_TL01_CLR1_char1_sprite_frame_control_frame_count_2, ZN => TL01_CLR1_n_11);
  TL01_CLR1_char1_sprite_frame_control_state_reg_0 : DFQD1BWP7T port map(CP => CTS_16, D => FE_PHN19_TL01_CLR1_char1_sprite_frame_control_new_state_0, Q => TL01_CLR1_char1_sprite_frame_control_state_0);
  TL01_CLR1_char1_sprite_frame_control_state_reg_1 : DFQD1BWP7T port map(CP => CTS_16, D => FE_PHN16_TL01_CLR1_char1_sprite_frame_control_new_state_1, Q => TL01_CLR1_char1_sprite_frame_control_state_1);
  TL01_CLR1_char2_sprite_frame_control_state_reg_0 : DFQD1BWP7T port map(CP => CTS_15, D => FE_PHN20_TL01_CLR1_char2_sprite_frame_control_new_state_0, Q => FE_PHN88_TL01_CLR1_char2_sprite_frame_control_state_0);
  TL01_CLR1_char2_sprite_frame_control_state_reg_1 : DFQD1BWP7T port map(CP => CTS_15, D => FE_PHN18_TL01_CLR1_char2_sprite_frame_control_new_state_1, Q => TL01_CLR1_char2_sprite_frame_control_state_1);
  TL01_CLR1_char2_sprite_frame_control_state_reg_2 : DFQD1BWP7T port map(CP => CTS_15, D => FE_PHN17_TL01_CLR1_char2_sprite_frame_control_new_state_2, Q => TL01_CLR1_char2_sprite_frame_control_state_2);
  TL01_CLR1_char1_sprite_frame_control_state_reg_2 : DFQD1BWP7T port map(CP => CTS_16, D => FE_PHN15_TL01_CLR1_char1_sprite_frame_control_new_state_2, Q => FE_PHN103_TL01_CLR1_char1_sprite_frame_control_state_2);
  TL01_CLR1_g1966 : INR2D1BWP7T port map(A1 => TL01_CLR1_n_1486, B1 => TL01_CLR1_n_1488, ZN => TL01_CLR1_n_6);
  TL01_CLR1_g1967 : INR2D1BWP7T port map(A1 => TL01_CLR1_n_1477, B1 => TL01_CLR1_n_1479, ZN => TL01_CLR1_n_5);
  TL01_CLR1_g1969 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_1487, B1 => FE_PHN111_TL01_CLR1_char1_sprite_frame_control_frame_count_2, ZN => TL01_CLR1_n_10);
  TL01_CLR1_g1970 : IND2D1BWP7T port map(A1 => TL01_CLR1_n_1478, B1 => TL01_CLR1_char2_sprite_frame_control_frame_count_2, ZN => TL01_CLR1_n_9);
  TL01_CLR1_g42007 : XNR2D1BWP7T port map(A1 => TL01_CLR1_n_517, A2 => TL01_CLR1_n_211, ZN => TL01_CLR1_n_1561);
  TL01_CLR1_g42008 : XNR2D1BWP7T port map(A1 => char1posy(1), A2 => char1posy(2), ZN => TL01_CLR1_n_1562);
  TL01_CLR1_g42009 : ND2D0BWP7T port map(A1 => hcountintern(8), A2 => hcountintern(9), ZN => TL01_CLR1_n_1563);
  TL01_CLR1_g42010 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_339, A2 => TL01_CLR1_n_1480, ZN => TL01_CLR1_n_1564);
  TL01_CLR1_g42011 : NR2D1BWP7T port map(A1 => TL01_CLR1_n_338, A2 => TL01_CLR1_n_1489, ZN => TL01_CLR1_n_1565);

end routed;
