configuration input_driver_behavioural_cfg of input_driver is
	for behavioural
		end for;
end configuration input_driver_behavioural_cfg ;
