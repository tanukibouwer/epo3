../../physics/jump_calculator_behaviour_cfg.vhd