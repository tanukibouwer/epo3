../../input/input_driver.vhd