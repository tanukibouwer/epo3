../../physics/physics_top.vhd