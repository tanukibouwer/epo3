configuration input_register_behavioural_cfg of input_register is
	for behavioural
		end for;
end configuration input_register_behavioural_cfg; 
