configuration Hsync_gen_cfg of Hsync_gen is
    for rtl
    end for;
end configuration Hsync_gen_cfg;