../../memory/m_writelogic_cfg.vhd