configuration damagecalculator-behavioural-cfg of damagecalculator is
	for behavioural
	end for;
end configuration damagecalculator-behavioural-cfg;
