configuration p_mux_behavioural_cfg of p_mux is
   for behavioural
   end for;
end p_mux_behavioural_cfg;
