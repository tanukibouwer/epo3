../../memory/m_toplevel_cfg.vhd