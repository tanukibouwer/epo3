library IEEE;
use IEEE.std_logic_1164.ALL;

entity p_dampener_tb is
end p_dampener_tb;

