../../VGA/VGA_frame_cnt_cfg.vhd