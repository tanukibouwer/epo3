configuration t_8bregs_cfg of t_8bregs is
    for rtl
    end for;
end configuration t_8bregs_cfg;