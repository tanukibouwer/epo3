configuration physics_adder_behaviour_cfg of physics_adder is
   for behaviour
   end for;
end physics_adder_behaviour_cfg;
