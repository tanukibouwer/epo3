configuration ram_8b_cfg of ram_8b is
    for behaviour
    end for;
 end ram_8b_cfg;