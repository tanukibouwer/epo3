../../memory/m_ram8bit_cfg.vhd