configuration t_4bregs_cfg of t_4bregs is
    for rtl
    end for;
end configuration t_4bregs_cfg;