configuration gravity_behaviour_cfg of gravity is
   for behaviour
   end for;
end gravity_behaviour_cfg;
