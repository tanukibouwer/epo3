../../VGA/VGA_char_sprites.vhd