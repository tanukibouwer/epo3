../../VGA/VGA_V_line_cnt_cfg.vhd