configuration H_pix_cnt_cfg of H_pix_cnt is
    for behavioural
    end for;
end configuration H_pix_cnt_cfg;