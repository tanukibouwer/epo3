../../physics/physics_system.vhd