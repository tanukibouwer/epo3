../../VGA/VGA_H_pix_cnt_cfg.vhd