../../physics/jump_calculator.vhd