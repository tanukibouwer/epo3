../../memory/m_ram9bit.vhd