../../VGA/VGA_graphics_card.vhd