library IEEE;
use IEEE.std_logic_1164.ALL;

entity physics_adder_tb is
end physics_adder_tb;

