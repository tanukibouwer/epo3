configuration Vsync_gen_cfg of vsync_gen is
    for rtl
    end for;
end configuration Vsync_gen_cfg;