library IEEE;
use IEEE.std_logic_1164.ALL;

entity p_impulse_add_tb is
end p_impulse_add_tb;

