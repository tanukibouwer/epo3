../../input/input_register.vhd