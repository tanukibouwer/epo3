configuration t_8bregs_perframe_cfg of t_8bregs_perframe is
    for rtl
    end for;
end configuration t_8bregs_perframe_cfg;