../../VGA/VGA_char_offset_adder_cfg.vhd