configuration ram_4b_cfg of ram_4b is
    for behaviour
    end for;
 end ram_4b_cfg;