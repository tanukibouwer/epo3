../../attack/coldet-behaviour-cfg.vhd