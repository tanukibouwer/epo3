configuration input_deserialiser_behavioural_cfg of input_deserialiser is
	for behavioural
		end for;
end configuration input_deserialiser_behavioural_cfg;
