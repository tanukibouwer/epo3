configuration killzonedetector_behavioural_cfg of killzonedetector is
	for behavioural
		end for;
end configuration killzondetector_behavioural_cfg;
