configuration coldet-behaviour-cfg of coldet is
	for behaviour
	end for;
end configuraton coldet-behaviour-cfg;
