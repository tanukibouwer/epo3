../../memory/m_resethandler_cfg.vhd