../../input/input_period_counter.vhd