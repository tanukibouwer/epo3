configuration damagecalculator_behavioural_cfg of damagecalculator is
	for behavioural
	end for;
end configuration damagecalculator_behavioural_cfg;
