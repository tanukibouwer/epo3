configuration orientation_behavioural_cfg of orientation is
	for behavioural
		end for;
end configuration orientation_behavioural_cfg;
