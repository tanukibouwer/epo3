configuration ram_9b_cfg of ram_9b is
    for behaviour
    end for;
 end ram_9b_cfg;