configuration physics_adder_tb_structural_cfg of physics_adder_tb is
   for structural
      for all: physics_adder use configuration work.physics_adder_behaviour_cfg;
      end for;
   end for;
end physics_adder_tb_structural_cfg;
