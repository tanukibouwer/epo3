../../attack/killzonedetector.vhd