../../VGA/VGA_number_sprite_cfg.vhd