configuration char_animation_fsm_cfg of char_animation_fsm is
    for behavioural
    end for;
end configuration char_animation_fsm_cfg;