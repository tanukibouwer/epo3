../../physics/position_adder.vhd