../../main/toplevel.vhd