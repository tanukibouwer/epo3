../../VGA/VGA_V_line_cnt.vhd