configuration orientation-behavioural-cfg of orientation is
	for behavioural
		end for;
end configuration orientation-behavioural-cfg;
