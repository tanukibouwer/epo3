../../physics/physics_system_behaviour_cfg.vhd