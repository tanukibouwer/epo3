configuration h_player_movement_behaviour_cfg of h_player_movement is
   for behaviour
   end for;
end h_player_movement_behaviour_cfg;
