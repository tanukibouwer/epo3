configuration m_resethandler_structural_cfg of m_resethandler is
   for structural
   end for;
end m_resethandler_structural_cfg;