../../attack/orientation.vhd