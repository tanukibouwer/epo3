../../attack/damagecalculator.vhd