../../physics/p_knockback_calculator_behaviour_cfg.vhd