../../physics/p_mux.vhd