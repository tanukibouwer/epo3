configuration char_offset_adder_cfg of char_offset_adder is
    for computational
    end for;
end configuration char_offset_adder_cfg;