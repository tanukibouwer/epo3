configuration input_buffer_behavioural_cfg of input_buffer is
	for behavioural
	end for;
end configuration input_buffer_behavioural_cfg;
