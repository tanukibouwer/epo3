../../attack/attackpressed.vhd