configuration attackpressed-behavioural-cfg of attackpressed is
	for behavioural
		end for;
end configuration attackpressed-behavioural-cfg;
