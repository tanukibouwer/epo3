configuration input_period_counter_behavioural_cfg of input_period_counter is
	for behavioural
		end for;
end configuration input_period_counter_behavioural_cfg;
