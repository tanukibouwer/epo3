../../input/input_buffer.vhd