../../physics/h_player_movement.vhd