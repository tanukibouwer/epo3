../../input/input_toplevel_structural_cfg.vhd