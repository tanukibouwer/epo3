configuration frame_cnt_cfg of frame_cnt is
    for behavioural
    end for;
end configuration frame_cnt_cfg;