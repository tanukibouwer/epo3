--module: number_sprite
--version: a2.0
--author: Parama Fawwaz & Kevin Vermaat
--------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------
--MODULE DESCRIPTION
--! This module is the static ROM for the sprites regarding the numbers that can be shown on screen
--! 
--! The resolution of the sprites is 9 x 20 which will be scaled up by 4 on the actual screen. 
--! This will be done by the coloring module
--! 
--! TODO: update this to become 16 lines instead of 20
--! 
--------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity number_sprite is
    port (
        -- clk         : in std_logic;
        number : in std_logic_vector(3 downto 0); -- 9 (max is 1001 in binary)

        line1  : out std_logic_vector(15 downto 0);
        line2  : out std_logic_vector(15 downto 0);
        line3  : out std_logic_vector(15 downto 0);
        line4  : out std_logic_vector(15 downto 0);
        line5  : out std_logic_vector(15 downto 0);
        line6  : out std_logic_vector(15 downto 0);
        line7  : out std_logic_vector(15 downto 0);
        line8  : out std_logic_vector(15 downto 0);
        line9  : out std_logic_vector(15 downto 0);
        line10 : out std_logic_vector(15 downto 0);
        line11 : out std_logic_vector(15 downto 0);
        line12 : out std_logic_vector(15 downto 0);
        line13 : out std_logic_vector(15 downto 0);
        line14 : out std_logic_vector(15 downto 0);
        line15 : out std_logic_vector(15 downto 0);
        line16 : out std_logic_vector(15 downto 0);
        line17 : out std_logic_vector(15 downto 0);
        line18 : out std_logic_vector(15 downto 0);
        line19 : out std_logic_vector(15 downto 0);
        line20 : out std_logic_vector(15 downto 0);
        line21 : out std_logic_vector(15 downto 0);
        line22 : out std_logic_vector(15 downto 0);
        line23 : out std_logic_vector(15 downto 0);
        line24 : out std_logic_vector(15 downto 0)


    );
end number_sprite;

architecture behavioural of number_sprite is
begin
    process (number) --inverted colored numbers! 
    begin

        case number is
            when "0000" => -- zero
                line1  <= "0000000000000000";
                line2  <= "0111111111111110";
                line3  <= "0100000000001110";
                line4  <= "0100000000001110";
                line5  <= "0100000000001110";
                line6  <= "0100000000001110";
                line7  <= "0100000000001110";
                line8  <= "0100000000001110";
                line9  <= "0100000000001110";
                line10 <= "0100000000001110";
                line11 <= "0100000000001110";
                line12 <= "0100000000001110";
                line13 <= "0100000000001110";
                line14 <= "0100000000001110";
                line15 <= "0100000000001110";
                line16 <= "0100000000001110";
                line17 <= "0100000000001110";
                line18 <= "0100000000001110";
                line19 <= "0100000000001110";
                line20 <= "0100000000001110";
                line21 <= "0100000000001110";
                line22 <= "0100000000001110";
                line23 <= "0111111111111110";
                line24 <= "0000000000000000";
 
            when "0001" => -- one
                line1  <= "0000000000000000";
                line2  <= "0000000000001110";
                line3  <= "0000000000111110";
                line4  <= "0000000111001110";
                line5  <= "0000011000001110";
                line6  <= "0011100000001110";
                line7  <= "0000000000001110";
                line8  <= "0000000000001110";
                line9  <= "0000000000001110";
                line10 <= "0000000000001110";
                line11 <= "0000000000001110";
                line12 <= "0000000000001110";
                line13 <= "0000000000001110";
                line14 <= "0000000000001110";
                line15 <= "0000000000001110";
                line16 <= "0000000000001110";
                line17 <= "0000000000001110";
                line18 <= "0000000000001110";
                line19 <= "0000000000001110";
                line20 <= "0000000000001110";
                line21 <= "0000000000001110";
                line22 <= "0000000000001110";
                line23 <= "0000000000001110";
                line24 <= "0000000000000000";
            when "0010" => -- two
                line1  <= "0000000000000000";
                line2  <= "0000111111111000";
                line3  <= "0001100000001100";
                line4  <= "0110000000000110";
                line5  <= "0110000000000110";
                line6  <= "0000000000000110";
                line7  <= "0000000000000110";
                line8  <= "0000000000000110";
                line9  <= "0000000000000110";
                line10 <= "0000000000000110";
                line11 <= "0000000000001100";
                line12 <= "0000000000011000";
                line13 <= "0000000000100000";
                line14 <= "0000000001000000";
                line15 <= "0000000010000000";
                line16 <= "0000000100000000";
                line17 <= "0000001000000000";
                line18 <= "0000010000000000";
                line19 <= "0000100000000000";
                line20 <= "0001000000000000";
                line21 <= "0010000000000000";
                line22 <= "0010000000000000";
                line23 <= "0111111111111110";
                line24 <= "0000000000000000";
            when "0011" => -- three
                line1  <= "0000000000000000";
                line2  <= "0111111111111100";
                line3  <= "0000000000001110";
                line4  <= "0000000000001110";
                line5  <= "0000000000001110";
                line6  <= "0000000000001110";
                line7  <= "0000000000001110";
                line8  <= "0000000000001110";
                line9  <= "0000000000001110";
                line10 <= "0000000000001110";
                line11 <= "0000000000001110";
                line12 <= "0111111111111100";
                line13 <= "0000000000001110";
                line14 <= "0000000000001110";
                line15 <= "0000000000001110";
                line16 <= "0000000000001110";
                line17 <= "0000000000001110";
                line18 <= "0000000000001110";
                line19 <= "0000000000001110";
                line20 <= "0000000000001110";
                line21 <= "0000000000001110";
                line22 <= "0000000000001110";
                line23 <= "0111111111111100";
                line24 <= "0000000000000000";
            when "0100" => -- four
                line1  <= "0000000000000000";
                line2  <= "0100000000001110";
                line3  <= "0100000000001110";
                line4  <= "0100000000001110";
                line5  <= "0100000000001110";
                line6  <= "0100000000001110";
                line7  <= "0100000000001110";
                line8  <= "0100000000001110";
                line9  <= "0100000000001110";
                line10 <= "0100000000001110";
                line11 <= "0111111111111110";
                line12 <= "0000000000001110";
                line13 <= "0000000000001110";
                line14 <= "0000000000001110";
                line15 <= "0000000000001110";
                line16 <= "0000000000001110";
                line17 <= "0000000000001110";
                line18 <= "0000000000001110";
                line19 <= "0000000000001110";
                line20 <= "0000000000001110";
                line21 <= "0000000000001110";
                line22 <= "0000000000001110";
                line23 <= "0000000000001110";
                line24 <= "0000000000000000";
            when "0101" => -- five
                line1  <= "0000000000000000";
                line2  <= "0011111111111110";
                line3  <= "0100000000000000";
                line4  <= "0100000000000000";
                line5  <= "0100000000000000";
                line6  <= "0100000000000000";
                line7  <= "0100000000000000";
                line8  <= "0100000000000000";
                line9  <= "0100000000000000";
                line10 <= "0100000000000000";
                line11 <= "0100000000000000";
                line12 <= "0011111111111100";
                line13 <= "0000000000001110";
                line14 <= "0000000000001110";
                line15 <= "0000000000001110";
                line16 <= "0000000000001110";
                line17 <= "0000000000001110";
                line18 <= "0000000000001110";
                line19 <= "0000000000001110";
                line20 <= "0000000000001110";
                line21 <= "0000000000001110";
                line22 <= "0000000000001110";
                line23 <= "0111111111111100";
                line24 <= "0000000000000000";
            when "0110" => -- six
                line1  <= "0000000000000000";
                line2  <= "0000111111111100";
                line3  <= "0001100000000000";
                line4  <= "0011000000000000";
                line5  <= "0110000000000000";
                line6  <= "0110000000000000";
                line7  <= "0110000000000000";
                line8  <= "0110000000000000";
                line9  <= "0110000000000000";
                line10 <= "0110000000000000";
                line11 <= "0110000000000000";
                line12 <= "0011111111111100";
                line13 <= "0110000000001110";
                line14 <= "0110000000001110";
                line15 <= "0110000000001110";
                line16 <= "0110000000001110";
                line17 <= "0110000000001110";
                line18 <= "0110000000001110";
                line19 <= "0110000000001110";
                line20 <= "0110000000001110";
                line21 <= "0110000000001110";
                line22 <= "0110000000001110";
                line23 <= "0011111111111100";
                line24 <= "0000000000000000";
            when "0111" => -- seven
                line1  <= "0000000000000000";
                line2  <= "0111111111111110";
                line3  <= "0000000000111110";
                line4  <= "0000000000001110";
                line5  <= "0000000000001110";
                line6  <= "0000000000001110";
                line7  <= "0000000000001110";
                line8  <= "0000000000001110";
                line9  <= "0000000000001110";
                line10 <= "0000000000001110";
                line11 <= "0000000000001110";
                line12 <= "0000001111111110";
                line13 <= "0000000000001110";
                line14 <= "0000000000001110";
                line15 <= "0000000000001110";
                line16 <= "0000000000001110";
                line17 <= "0000000000001110";
                line18 <= "0000000000001110";
                line19 <= "0000000000001110";
                line20 <= "0000000000001110";
                line21 <= "0000000000001110";
                line22 <= "0000000000001110";
                line23 <= "0000000000001110";
                line24 <= "0000000000000000";
            when "1000" => -- eight
                line1  <= "0000000000000000";
                line2  <= "0111111111111110";
                line3  <= "0100000000001110";
                line4  <= "0100000000001110";
                line5  <= "0100000000001110";
                line6  <= "0100000000001110";
                line7  <= "0100000000001110";
                line8  <= "0100000000001110";
                line9  <= "0100000000001110";
                line10 <= "0100000000001110";
                line11 <= "0100000000001110";
                line12 <= "0111111111111110";
                line13 <= "0111111111111110";
                line14 <= "0100000000001110";
                line15 <= "0100000000001110";
                line16 <= "0100000000001110";
                line17 <= "0100000000001110";
                line18 <= "0100000000001110";
                line19 <= "0100000000001110";
                line20 <= "0100000000001110";
                line21 <= "0100000000001110";
                line22 <= "0100000000001110";
                line23 <= "0111111111111110";
                line24 <= "0000000000000000";
            when "1001" => -- nine
                line1  <= "0000000000000000";
                line2  <= "0111111111111110";
                line3  <= "0100000000001110";
                line4  <= "0100000000001110";
                line5  <= "0100000000001110";
                line6  <= "0100000000001110";
                line7  <= "0100000000001110";
                line8  <= "0100000000001110";
                line9  <= "0100000000001110";
                line10 <= "0100000000001110";
                line11 <= "0100000000001110";
                line12 <= "0111111111111110";
                line13 <= "0111111111111110";
                line14 <= "0000000000001110";
                line15 <= "0000000000001110";
                line16 <= "0000000000001110";
                line17 <= "0000000000001110";
                line18 <= "0000000000001110";
                line19 <= "0000000000001110";
                line20 <= "0000000000001110";
                line21 <= "0000000000001110";
                line22 <= "0000000000001110";
                line23 <= "0111111111111110";
                line24 <= "0000000000000000";
            when others =>
                null;
        end case;

    end process;

end behavioural;