../../VGA/VGA_Hsync_gen_cfg.vhd