configuration killzonedetector-behavioural-cfg of killzonedetector is
	for behavioural
		end for;
end configuration killzondetector-behavioural-cfg;
