../../memory/m_ram4bit.vhd