../../VGA/VGA_screen_scan.vhd