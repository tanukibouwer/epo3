../../VGA/VGA_char_animation_fsm.vhd