../../memory/m_ram10bit_cfg.vhd