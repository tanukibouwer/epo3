../../VGA/VGA_char_sprites_cfg.vhd