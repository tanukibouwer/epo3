../../physics/velocity_interpolator_behaviour_cfg.vhd