configuration jump_calculator_behaviour_cfg of jump_calculator is
   for behaviour
   end for;
end jump_calculator_behaviour_cfg;
