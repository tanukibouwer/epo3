../../memory/m_ram8bit.vhd