configuration h_pix_cnt_cfg of h_pix_cnt is
    for behavioural
    end for;
end configuration h_pix_cnt_cfg;