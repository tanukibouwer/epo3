../../input/input_buffer_behavioural_cfg.vhd