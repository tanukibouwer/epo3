../../VGA/VGA_frame_cnt.vhd