../../memory/m_ram9bit_cfg.vhd