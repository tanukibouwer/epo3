../../physics/collision_resolver_behaviour_cfg.vhd