../../input/input_deserializer.vhd