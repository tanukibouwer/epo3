configuration killzonedetector_behavioural_cfg of killzonedetector is
	for behavioural
		end for;
end configuration killzonedetector_behavioural_cfg;
