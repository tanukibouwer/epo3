../../memory/m_writelogic.vhd