../../input/input_jump.vhd