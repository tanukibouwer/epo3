configuration ram_10b_cfg of ram_10b is
    for behaviour
    end for;
 end ram_10b_cfg;