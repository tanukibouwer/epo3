configuration writelogic_cfg of writelogic is
    for behaviour
    end for;
 end writelogic_cfg;