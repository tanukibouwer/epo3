../../physics/gravity.vhd