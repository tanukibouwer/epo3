../../attack/toplevelattack.vhd