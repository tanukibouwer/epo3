configuration V_line_cnt_cfg of V_line_cnt is
    for behavioural
    end for;
end configuration V_line_cnt_cfg;