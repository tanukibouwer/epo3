../../attack/killzonedetector-behavioural-cfg.vhd