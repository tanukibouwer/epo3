../../VGA/VGA_screen_scan_cfg.vhd