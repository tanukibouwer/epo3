--module: number_sprite
--version: a2.0.7
--author: Parama Fawwaz & Kevin Vermaat
--------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------
--MODULE DESCRIPTION
-- This module is the static ROM for the sprites regarding the numbers that can be shown on screen
-- 
-- This will be a modular component with an enable signal that will allow for the component to take over
-- coloring duties
-- 
--------------------------------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity number_sprite is
    port (
        -- which number to display
        number : in std_logic_vector(3 downto 0); -- 9 (max is 1001 in binary)
        -- data to go through the array
        hcount : in std_logic_vector(9 downto 0);
        vcount : in std_logic_vector(9 downto 0);
        boundx : in std_logic_vector(9 downto 0);
        boundy : in std_logic_vector(9 downto 0);

        R_data : out std_logic_vector(3 downto 0);
        G_data : out std_logic_vector(3 downto 0);
        B_data : out std_logic_vector(3 downto 0)

    );
end number_sprite;

architecture behavioural of number_sprite is

    -- integer values for the counts
    -- signal int_hcount, int_vcount : integer;
    -- signal int_boundx, int_boundy : integer;

    -- declare the array for the colours
    subtype color_val is std_logic_vector(11 downto 0); -- R(11,10,9,8) G(7,6,5,4) B(3,2,1,0)
    type num_sprite_x is array (0 to 15) of color_val;
    type num_sprite_y is array (0 to 23) of num_sprite_x;

    -- fill the arrays
    constant zero : num_sprite_y := 
    ( 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")) 
    ); 
    
    
    constant one : num_sprite_y := 
    ( 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")) 
    ); 
    
    
    constant two : num_sprite_y :=
    ( 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")) 
    ); 
    
     
    constant three : num_sprite_y :=
    ( 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")) 
    ); 
    
     
    constant four : num_sprite_y := 
    ( 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")) 
    ); 
    
    
    constant five : num_sprite_y :=
    ( 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")) 
    ); 
    
    
    constant six : num_sprite_y := 
    ( 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")) 
    ); 
    
    
    constant seven : num_sprite_y := 
    ( 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")) 
    ); 
    
    
    constant eight : num_sprite_y := 
    ( 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")) 
    ); 
    
    
    constant nine : num_sprite_y :=
    ( 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("000100010001"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")), 
    (("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111"),("111111111111")) 
    ); 
    
    
    
begin
    -- int_hcount <= to_integer(unsigned(hcount));
    -- int_vcount <= to_integer(unsigned(vcount));
    -- int_boundx <= to_integer(unsigned(boundx));
    -- int_boundy <= to_integer(unsigned(boundy));

    process (number, hcount, vcount)
        variable int_hcount : integer;
        variable int_vcount : integer;
        variable int_boundx : integer;
        variable int_boundy : integer;
        
    begin
        int_hcount := to_integer(unsigned(hcount));
        int_vcount := to_integer(unsigned(vcount));
        int_boundx := to_integer(unsigned(boundx));
        int_boundy := to_integer(unsigned(boundy));
        case number is
            when "0000" => -- zero
                R_data <= zero(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(11 downto 8);
                G_data <= zero(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(7 downto 4);
                B_data <= zero(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(3 downto 0);
            when "0001" => -- one
                R_data <= one(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(11 downto 8);
                G_data <= one(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(7 downto 4);
                B_data <= one(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(3 downto 0);
            when "0010" => -- two
                R_data <= two(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(11 downto 8);
                G_data <= two(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(7 downto 4);
                B_data <= two(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(3 downto 0);
            when "0011" => -- three
                R_data <= three(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(11 downto 8);
                G_data <= three(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(7 downto 4);
                B_data <= three(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(3 downto 0);
            when "0100" => -- four
                R_data <= four(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(11 downto 8);
                G_data <= four(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(7 downto 4);
                B_data <= four(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(3 downto 0);
            when "0101" => -- five
                R_data <= five(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(11 downto 8);
                G_data <= five(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(7 downto 4);
                B_data <= five(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(3 downto 0);
            when "0110" => -- six
                R_data <= six(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(11 downto 8);
                G_data <= six(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(7 downto 4);
                B_data <= six(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(3 downto 0);
            when "0111" => -- seven
                R_data <= seven(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(11 downto 8);
                G_data <= seven(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(7 downto 4);
                B_data <= seven(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(3 downto 0);
            when "1000" => -- eight
                R_data <= eight(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(11 downto 8);
                G_data <= eight(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(7 downto 4);
                B_data <= eight(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(3 downto 0);
            when "1001" => -- nine
                R_data <= nine(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(11 downto 8);
                G_data <= nine(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(7 downto 4);
                B_data <= nine(int_vcount - (int_boundy + 1))(int_hcount - (int_boundx + 1))(3 downto 0);
        
            when others => -- fallback for error handling and checking
                R_data <= "0000";
                G_data <= "0000";
                B_data <= "0000";
        end case;
    end process;

end behavioural;