../../memory/m_toplevel.vhd