configuration input_jump_behavioural_cfg of input_jump is
	for behavioural
		end for;
end configuration input_jump_behavioural_cfg ;
