../../VGA/VGA_H_pix_cnt.vhd