configuration dig3_num_splitter_cfg of dig3_num_splitter is
    for behavioural
    end for;
end configuration dig3_num_splitter_cfg;