../../input/input_deserializer_behavioural_cfg.vhd