../../attack/coldet.vhd